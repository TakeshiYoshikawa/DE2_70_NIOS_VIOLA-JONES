��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�oBy��hk;��k�X G���2��LO���N�=�qs�W|}���O����9x�IN(^�?�@�\����Dם��ُ�|�f(��F����Q�V�ӈ��1��'7#w���C�Pn�+�|<	 �f�����L��
���i����t�p����Ppv����^M��TV��I��6�.��L�Qf�*��
`�<z^0�^�����q:Ѿ��!�y}��`���@��u'y��j��,3!
cI��2jp�VX��/���C���Q��JI0BT��C��㛝����
'r �%�/�|p��L:o��:��v��-����볕­�(�u
U��,�Ƃ���(:;m?�|��`E�S�T�9�_��i��~�lܴqzx��&�N��bOYw�iTɇ����16��i&C��T������4	����K�Р4�A|���	��x�c;�;�5�g�������[{T�Ro�J�j��Γi��&��#.D��5��龥w�0V�"���F�!gԈ�	�������0�¥(�~GR8�&~���ä\��"�u���ٱ�?�T�4���A�T�.�������E�$����,\B�F%�j)�%eb�tm��?�[�e]!_Iz�)�x���1���Z��d,M��U�	�ݶY��o��+-����c 2Ǹ���������V��B�}�#�����]��q>V�h����M�����_��kۈ�sax�0+N}"M(�Xw/��l�Ů'm�1uP�
̜���nːtߐ{��L��IkC�
�ʏ*)+��7ӫ4�瑄���򾝯�c
qe��,O1�c曧��B�)Q���[��j��L�N:���Z'7�W�i��mz������.;NF�2O(F龒"yOt�?���D�^�ad�/4�ޑ���ɰ��˹\2�Э�i�ط#3,W�	�q��e�,�T��]�E�E�^��iu��)��@&���"��Q۽?����@ ���Jq(������b��xk��6�Lx��E9M���" �c\�bh�?C���(9��탁�.[�{��G��H�:Q�%��sh��V0%��$�W�wQo�v�6;�Î������	�|�{�����ϩZ��q
F�4P�L�O����r�M�.T��x+�M��{0��r��&~�6�iѦ�uNԦ��jV�fb��@��eiI�R����j�:�9%֮*Ϲw���K�bFQg_��A)^w\N姖h�L�C�����f���L�5��OM3eB3[�H�N-$���=�^�t(_�vi%/F��ׯX��L#.*o�^�2i�@�M���d�˶�KQGف�8�y�U1�ۨ��P�ӥ��aE�Q!�8�ӻ�ԉ3-���}�2B�-��/Tqp��hQ�I���o� ]r\h3��M�Nf�M��5���ݘ*�>���l� �u�Ol����e]�Kq��q��GS���kAR;8ef�]��!�<l�ƈN2as��r<���ym�]�G��R�s5	G�sd�V@���[�$MA����iȼ���j*�_�271yy@�0�o�Փ�*ƇO��Q@� ��&?����1vo,���K:�����]�����k�,�4��t���R* Y�H�.@j�NM� ��'��|R���֫��a����U�
CNg���h��x��C4��.�WK#��td/^�Ja�������~�Msު�{+��m�i�\��E��� G�<C���᧸o_���D=4�~}�Q�+]#~4����,�ÿ���3���O]z����!{x=��/����1$zr���e������o���Q���|L)��E�lyzv�`���"K!�R7�$#^����;�vVFy$+9C1M��W[��5�d�8*K\w c����j2��ڋ��1d��זN�7�c�:0��%�
_�wMb6��)o���9�kɲ�O������K:5jv�����tO���*R%�X�{����[\�-=&k8xtώ����A�#��f���MX��xYvPn��D��!i .��2�(}l�\��G���!���Gj��RH�ݣƹ��w��wV�x=�\�U� ��bY�)%���/\���P;��FE���Nancz�@�(Y�7��1�x�hb1ձt��f�D^����:{[ڨP�H�ln���(��hWU���\�5U�ܗ���x"���p���I 臸�X<�{[�V��1!��ڛ~A*=�g�vGhT*{-�K�S���0�ԓ1�?1I*��B��v�޳�տ��4�>WCg�ÛJ
7�������·\�]jɞ�-�ė�N�7B�zQ�b�P����:�=2��'�5�Qq��n�D��X�xq�?*3䀃,��48NH[�c�r[���n���x+�Ɖ��eU�/?(�y�"5��G�,2�zMo��)�ٰy���V�j���1���
�ÔʒX�f�d��P[�jGϞ���m�^���0�f���g^4y�hH�l�2�fI���}�I��]sU~��L=T:����]�}��C�׸+WZ�'�{q�����O� 8L.���z����;P����m~�
|F�ÙM�&���h��sG�Yc������2d]t�X��V��Ϙ�´���i�^�t٠���< re����GF���b�"��=��W��t{(d0���!D���2���M�"n�X�� ���`����O������=Mc������E�bbߍ�v���7
�xė H5�&�Hgcm٤4h��6�6Z��a(� �)���{\�4킵�z�΃%�3�ώ��&��k<i��:�&�C|G���s��ݨ�G�.��4�����'�����1x�����8]����K�&Hj��,ͣ��MC��7a�u����IZ6F� ��`7��[�`���c�bC����8{��i�ka[P��e�/���M���!Jv��`��xVo�Q��#|��T�����	W�� ٠Z��9K��#���OD ��O�9^���̚&��CЄ�}a(W��:��
��{$��=�7F`���6���$���ӻ�+LzZ�Oy]~{���*��MVV%�u�c�a��R��d�	�;I,@����܊��n?JU�ݙ�ڷ����L=�Zf�\ɲ�w��;Om��I�Ų !�������4wS:���,�3�L����*@�dk�
IL���[(��̚E!�j�5qo���b�V��N�?��_�j�&��ˇ"vʌ�8|��!p�jq�rG��2�N���Y��k}a4���݈j��Ov�t�����-��'e��hҷ&����}_�/����󓼩��3� 䧅��[=��a����9F-����i=K��Y�c��ݵ̅r0���4��"'�6DP���
v>�&Y����ă��D�"��+��O``i�B5$���/F�__�n+]U �O�����G��XV�A>[[	�-UV�c�� ��1 �m	�v�Ҧ'���Dn9�u��ifC�.����*%i�7ε*������F�yt������g,t�v6j�<��P���kx�ߵT-���sa��Cz~��l�0���6���O�!�٤���.H��6�g��g'f@��P�u_��ªځ�)�_}h�	�Q�'K4���}�kF�~���	�c��ޝ�����d�~&�ŭ7�'�BmO��h�k�8-���ȏ�L?}r�h�(��y�~�W��*�����*h��۱�+p���K��v�n/Yj�g^*|3��V7M��ˌV���R?t�����W�]�u��T�����,�bE>�������
���7S���8"�Xh�%��^��kuGe�����װ#9���,RΆ�5�)�Lh��=|մ��G�H$N3'r)y}9��������w3�n�_�a$		���=㡴�/d�gL���
k�W���"a��
q�L%�UR���w<���H��]�x͟�
:��P����_�oSʠoL�;g�TuҷŁ�_�B��޿1���5�C�rZ��Ѧ��uj�9�76���A��`��M��Y3��r��Ilq�i��n�&nߎ���v�s���[ 0+��3�KM���f��l�D^{t� ��	O��i�ܪ�q9؛�Z̍ޠ��P#,��Y�k�W�S���#�<Pc:>��fƉ_�b����M�+���e�ށZM�>���A5�1�2KNظYn-���A``���>x�:N�K�A���5�#�����6"��/�!>��͟����7��+�*%͞o���<r���5$������8���2v>hi]w&p��w�� ���#�$�u4�6�h�Wk�&Z�=��!��Y�>0�I$P�U^�@`�C�|�:S�����sD���*N!�YCf-44���yI�����+�+Fq�L'�45�C| s'��=��q�����}��cU�&��aY���Hk��u������.OgߡDs7�����&E���Κ 0_^D���Gg�(��O�I̟���"��H@X�yd���J��I!�}�l9=���YS:�H�j<��WU1FS�,W�F�i����F�VD�`��b�ۙyǽ�"�5:�>���]�{w���!����BC�+�79|�����݌R����?	`+�O�^^1�&��t%������?v��8@�h�=Q�K�7z���_,��t�;MmB]�t��/JZw
�[2�\����0��BL�����ܷZar>G��&���Q��\,g�f]p����%z�q,i1��?G>"�dw���ۙ��;ts����?��p�zr��d��+�y������$/�������l!��M`;�ذ��2�@&wFp�����m8�@4�ۮ/\e�G5-�Ll�	�}we�bB�U�s#<p�Y�@ٸg����5�'�ʌ^q��g�p���6$x��ԩM8���ȸ�����	�������R''��A� o�?<f�����D�ш�$&C<�V�[V��h!�� �8�+��\�Џ�56����˰��0\��5������{W�䨈Vh0/��F��modvF~<��X�pV�E�?jAE7-ԣ�p�����Z��Qg����x�D�+v�L���b��nC͌�ꌈ�J�[[��=R��`�)2!نJwAX@���#D�4L���|c�LT)�P�I�)��5Ex��`��7����`qv;��?,!I���@'�H������A$�Ԋ�c��v�5�\��H>�P��Μ+�|�C���.�ˑ�չu�E�;�X�YHE\��w�'qT�	22l�-ǭx} �R9��|�W N�&�}]t}��jS��#�M�t�u�W����G�qQ�E�&6�,��Ry{�Sv/��v�>K��ES�%��ط3P�X���|��?G�WR|�������`/`{�gV�c����G7����lB���ˏ��	����ݚVY�+C畱��]-tp�s��g��U[_gg�ߞ�<� 4��1^�agY�c���U��Ǣ��^�����_!��ڸ�ZW�����zq��W}s�t�uD�eT�X�P51���ţ9��Y��ڇk7�^��!��#7�d��&�q���g˚�do\��f�u�Fc]8�úF%\���K+m���.��ܣn��ʱ�D3 uĕ�3*�*-�\��*�I�Yp�IV��솳B�hx5`aLn�S���[J�T]�@C-���݆y�;��	�F����¬���w��F��|%_48\��̫K��A*��ڨ�
�`%��b��'�6nl(�S����k�0:���L����r���qptd�����2k���j��|!�V��~����s�_���@>���"��ݞg2F1%���L��%��EI���wJv��Yۂ����tg��1+	�Sb������x��Tu��"i�҆x�G[0�����^����,BP�z��+֑�� M����@�e�?5�Z>jŸ��g�9,4*��+\f"�cP4�(3�-K[��96�ρt�%��7b�u�7�c��H����x%>o�0^�X��7���,��N��ﰑ\�	M{3�J)��oa36��gh�@�k��3u,�6���+�.�'���!�-��2�u��AfL����L�6��%�Pmv��/D��:�]��0�Eɱ���Iy�yW���@�܋Y��3�����v}�4x���N;���<]MJI����4:�'ω�
�H{����!y�Ċ�G�{fi�I�����dG��r�nʦTg%����Y�}��@S���L�+k����܈}<�� �,�r+�CͶ��w�q������7�7�����1�j[�ß�z����T�'L�3�w,H�D%������ �3�$�G铮K�k�3�]�OE���h���r���Yc$��QC��Z��˛�zY_n^���kļ3,~�j��Ǫ��dsR�JhW[�g�G�� �5� ����������w�'�����9O��05H)����=τ�в[{]��-,	o�	%ԅ)s~���G�(�(_(�9�DzaZ�K���=�5fj��O~�f��ҵ�,�~Oϓ{m��EY��@qq�L@"���|=�_Xo���A��l�H���C������0���D4+�Q )��arSq=�<�~3�����Q�st�q78x&�G�7t�B��ύ~�uޡ�����R���BIt�?N����4���J�4Jr(I�ص,6��^�(Ռ5K�T����">*)�y�?��׼����vM�uZ|kJ���X��(�j$�7�m�e����Npװ�	G�Q��>E���'; ��y��C)��h�`��ll���SwDkE죢!� ��=;�E0��#)`݋FFש��c�ҳ�5mIN����������n�j����[?H��n-ٰRXbr&�Ɇ���!��A�C�=v�f��B� �|�{9t̚B��/e�0z��9��Wn/�����ޭm�sB�q��ډ��%��%��G��f>?��v�y�ؗ���x�eQ�"��C��~lz����} =�^OH������W�(��e���L���'�O�A_�:�'cQ"��ħ�a�Z%���> T�p��2p)�PU*,����_s$t��(��S5(��:���v~�#6A�H��t�0^~�(?}�<�9����̳��-���X���1I�?5�� G�.�j ���/��������ӽl�qg�W�OBH�XE��A:Rh���m}8���Ƣ�k�\����s2K$tb�(6U�G.'��t�R��5���TM�������BP������¦U}i�p�L`w~ⳅ4�+�OY�#��w}U!�)�l��Q�۸*?%�b�ݳ�v��-<�� �����y+[��,��pȬ橵�%̇�q���E�2�8�6��h��p��B�OI��+�Xн��a��/![�
��:�����C�Rd���!��z���@��\�����O/�`�U��$��ܺ��#��5z>lȔ?b��kzh0�i�^�pݿ�`�m��6	��9yu����_:y9�C�6d�2�vg4�ap�eG}֔r�^H�G�Adrt;c:�TΨI���6��4����Y�¸#Et0Xq�g�^��(�|>�l)�U������x���q�JlFz8�<7�����N*h��
�n��sw����G|�c�]eAu�t��T8�E"|*K @A�?ޖ�;�s!'T�۱h�
�,1�xE~��psDLf���Z��;׈i3񒎮��ͬ&�H���id �B|��<��q.���%��,c�����ЯI	�fg5���������Θ��Q�.os�-��]	�#33�W#+d[����UV>��>��"̫4���R���q�G�G���qH��Ӈ����d��R��3f7���QU&u�q&�� �u�{��2���Z�>�!����"�@��j\�X�0!����5��� �H�<����⍐0"&�У�ٳD��/���t'&[�3*qD#�/D�i�>{�xS�)MiQ#F����u�ۅJ
���a]�e8��U/���2�E,;Zm����3�$�<i�R��êT�kBޣ���o�	dl��E> �/������ƶ�>�+J��ATA�UBʊ�j�Y�|"�����
�i�Q��"uj,:av"���ܳ����zg���G�����Dmecc(�Ю���^�:1!�ޣ!$��J�U1�f�-�Y�8H�|XH/�&}��Mպ��+<�_��F�^q fήK�I��:�Z��<��OO;VAJց���q����<�- ge�\��Ȱ��a(�33`f�E,�ɛ�w#knL~��ED�E�
��
��Jc,H�5�(���u���=.c�6�����+N��5���H͛hG&�'����t�d/-�.|'���*�@��DM������W�:f�>�;�f\ѕ	h���T�7zX��ep����Yt���ry�?�ET���<S���Nm��%�g�;;|�L8���S��E���������
��G7^��>h��R���@\5���]�����wt@��!!2��E�9�1_s g��͢])l��!^C�U�2�:W�
�Yc�Ϲ������v�Ȼ�Qɾ��4�ض U}�ٳۏZΆx�ᵳB�������	���vT	���'�`�d
�e�3R�~*��D�?
�~�^��f��+ð_�,f��3��d���,��fK�`���P�|�Vt�b�C�<�!�0�Xq=֙�➆��d���:A�U�.�aj��]~�I{�����_[%����?��g���{$����8߬�>%\8/�lx�"�Y���YMc\�~))��/��%`V�L� ���/��ֵ����N$��)��.1bt;�����l#�W�Sd�I(���2_tI�[�	M}�d��oY�&��nN�B9�?���7���� /(�j�Y�'Zqomqr0:(�U��"T��b1-�\���"��=�=�!�����-ab�H̯		��^r��v)v���1�/^R�����!;^WB(m���Օ4!WZ������[��u(J:}3UŲr������ �������5B�xs�]��2��M#�;c~.��_���St����i"��%
ܕ��]c�Mg����t�J��ݟZ�rk�$DN�
�t*b+����m��[x�n�h�J��`3o�&����Au{�
��(��nP���G��֞�Nak��a��u�PU�l��N�1zE#�B�D^f\y4
��0�b��_�6_63<���:@P�w�H�����N�H��Cַ���&I{ҵ�A���T�q/��Tˌqx�V�o�����q�v��� �{��L�to��������P�J1`�'�tn�H�s\u���Q�\���f�lr� �,�C-�=p0�L��YL��4:�r��g��{�� V/3��"D�[�f�ȍNd�zʭ�\� CCA����v	�e�m=	bYd�tD��pFZ3���*�͚��E9���*Z��4�(2A�}Y�����A0Ȟ��f�����m�9Z=��9Vm����^�^�;�"�^�cK�bJA~y96&ǆ�b^�!๋�ij{�������0;.;�q�!�i�\]�b�� )SL�`m'��:Yn�i���m��m?�����/�.���\($֧��*��߻?�;�Y8lxt��Q�EW���1ԩy\��`�i�eu�`4�ԟI���d�gu�W��g�^�O�i�:Bw�3+N�^��f��N\X�v�m�i
Ƴ�k�ֶDD梨I���
d���Q�/U�?��A�J�LD�;�P3�Q�s���>v��x�X-��n �o��n�'~�b��W���<�^Z�fY��2	p@���6�eJ�����IC���?�J��R范h���x�4�2��r����po9�ΧEn��-��V-���wS���>��*`Jn� ���$����J�_+�����s���v�gA�����9;�27p�X��.�
av�6�%�����_q]��5�C��I#k�`��i^RB��He��m�_�yWv�o #{I���n#-2A�,��tr���,�}	D�,���sY��c���`W�MC���"�
/�~q)V�/��K?1�g��J�|u/�B����d�.K�'��N��_�Q�`��@�Bt���M��8�[ �C�A^~"��Wwh�G�:0HŪ�/N���m`I+�f�8�ika
�p���
�j��59DZ�T���-�A���4�U��?��0B4]�:�3�/v�}"4[�WL&Q:�F��W��j�P�Lv�:�w�"���:��<���e>���T^�嘲`I:H�24���F?r�Z+?�{G/N�;�ӎ�0햂ݧ�:�1��j�Qw��ӿ}�W7�?͎ƜN��}�_jc-����;�^��Tsw���AS߹�g���@�s�yG�rWx��z�V^���2/e~��ٜx4�n>���p.0q\�V�=� �B@Q9�00>m{�K�I"+1�,�"�@�iV݀�Y�Sux&������z�	(��6BR�D��ִ� �EXg0�A�DBr�ص�)��f=[�ө�g�<2��������b�ӄ�����9�|˝��rI�}<��璊�H� ���ʗƣ����8V>n�	ƞ:�_Z�B���G�J��^�k���
C�c^-r3��ax�G��H=�)�Ϯ?�2��k��:��=�_�C�EK,>	O9��|�Ê"~��yP�O��U��Їx�u���r�QޕZ�y+'�W�x��5}(=W�6 ;cdx���nehk�g�2q>x9I���[vS#�������H�A���r���	���Y��:�ڌH�ML''.��K������i#��%�
���oϜH-�����{o">���+��(r�df�S����-�]LȮvc"�Ԏ3��>��� d��)��Kq$u5�FS#,n���=��f���+I��\��Y�]�(Oږ�*ģ�,��'A)E=����IH
��Ϻ!��v��0"_��mP�����V���-c�T�aG;_��<_a����b�P"��L#'�L������.�P��zt!���;�ibi��j�l����9�DҸFf[�X�O7*���B�^�Y������'U^֍�@�Js�)��ЉX�̭0m2B�R�a��w�F�jo$g(�V����øko8�=�1˄��U�B9VR�r�&o8-"�uw� �VZ��S2�=I�Z��﫧�5۫��(�Q �8}O��Y�ք�8`�Nz�<�X�/<�& �BR��֦�!�3�����hގݳ�zRI ���df�}��u����t@h&-�L\b�܆���;�e��iS��K8��2ĜU4��~�����HI����^0�!d!O�{Ɏ�`b��4��z�>�_%���Dr!M`7������;�/~���S����ik(�j��7!�;�2b�r-4��I�%�׀�Up�s�V��������?�Bs�/��A��jiqj����ڵ#P*)SR{å�h��-dnX�ɎG���r���TsY�7C��.`��Nz6�]4�q�5H8fh��tO���Xd��w6_��)D���|l��q���(2��@���G����*�ei���3R��tY����\��͎n*;��;�T
�<�
��b���|]d�5n|�^�me�wq�1�0�U/�)��Y�	�S�͐׺���]�]U��N�0�w��X�_���ѧ�k�	���-�8��~�!�]�.�߱Vur���S�(��;�ES�V0���>�u�'��{-���Ω�����2����z���&�h'�<;��W��r%��崵�6O"]����nT_pJbW���n����q;��g)�۴�RnX\Wi��z.��"��
�+
�i�Mi¥�n����\���8�U��vO�ɲ�:x�=�@��Ǯ����pt�mɴv�&��_�����0����c�fɱh�1�"�حƺC��\� ���n*�)ĝ����W��F;B�!.��V��J2�b�ծ���훏��@��W!��e�o����}Ѕ��L��s��<5���B9�_��8W�RGZ>��*x2��4&��u�$�};�*��7�1M��I!|�Y�Ɛ��6M�"�"\G��k`ļ`��c�y�+`?�΂2��Y�m�����_U�=�k�o�'�P������
�H���A4�W������3:
|>3����a�vq�jH��z�i�}�3�p1]P�m\T�B��1����4��	>���knt������IB6n+j�;H��O}ہ��g7��k*��Q��PD�#�� �w�q�v�JU�������&��|
>˫��q��f~���]g	Cn��j��Q��6�eT�,���+����"<�6I%9bxj�(�k���§�0\�K�Q�qdH�aVW��A@������'v=�ћt�����.�����xU�"��A�t�XO0�/A1��ХXi^t3�B#��~D�����gڽ#@���Z[!K�xdkٵ'�dA�}��L/��[�Ɉ��j���A`*Lw�t�	�%��u�i��c�mE'}"{3�/�2�(H"9�J!��[���!ˋ-��
	��%J����Ὦhou3��@5PR��D�N�/�0��Fi���l�jPN�MD��`�@6�]6�Zm8t�ؖC�ȏm����q�JB��A�i,��������PI���Zw7��p��U�/J'%���FC�L0X����]�<���#tk�a�Ѐ7����)r�k#�r:�XKY-�21��5z���q5��Nc�Q��_��]��~�)׫��\w����?��r�����hb��Ǖ�I�� �I��5�v$��^����T6�)���!{֢�U�F�j\E!1PLX,�2_��bsLE<���O��gJ�:�%�o�����'t�#:���Ҟđ��ŧ���!�8=I�*���+�cT��t��,X�G@xC���{sQ����Ae��!;���ʍ�fx9��]��hD�V�:�-��k �O�O�}��BpY!W�yb�������}�f4�NB��K|W#P�2h6jAg�R�Ee0��
���N��#L�Z.�\ME��D�ɲ3��;����K�Q�\��X�x��eǾ1VއM،v�OF����˟U����ۈ�k^�����n���6��Hht%�[�
��m��.�%���mӃ5�k�l�h\�%�5�\� ���Z٘��E��`,�~]/�EO��!��8��VnϋS��y��]�����I����9��>�Y�E�a��C\���,�,�OD��l�S���f�Β{�%�)�`cX�#du��Zd��;"�U���o,�88�%�Ͽ�M��52���]	�*:����G��C���M�i��+g@�`J��d^�J�H����u� M*�H[OR������gZ���[{�Z�*�(�@�>x�>,�:<����<����zQ��#���V���4<s@((A���k��d���Th��@�-:U�{h�g��݌q�.��te���i��e,g��<[���gB����:%~���g�@RT��l�Q4W�# |V�gNl<���\#�� ��D5	���ô� \�
��Y��<���,\5����1���>�a4Z%�1c�&�����}X�m��	d_�~�y$�1uN�ud�(�Y����j�C��Q	�y��/k5	_�3�w3.y��Yߛ���� �rJF���f��sk�`ܽD���9�{�Y S���nn����M�S�er(��|�=M��{4��(v�A�$WT��`7�~�qd�c-=2�'ѻ���~6v%�$(8��5�,����� �/҈�:6�8�*�.#%^�y�r�z?bkǇg��G;�=�YM�����kE���N�(5���c���
�r����6��>�7�T�3�>�v�5Y兀����>U#�o��$ Gj��
�Y;^���&@˩�4^�N�6��_�Ǻd	 6UD8�YnD��S8I\�-�,��=LD��/N)���\�B��M�Zp���f�	2բ���VM�şf��ĉ�ʣ7���}B����O<�*�n�):_�"�`�	���~ߐ)��������w��Ć�g´B���mr����蘉F�D��j�a��mc`�?hKr��[�,�#�R�5Mw�W @3|�>��uq��M��,������Y8DT;3,��a�1=zf�VA��[8��U�J�MA���3Gg�w;�F҇���8�6��[4�n8���˘�~���G�^�Qt��������(�v�BC�����q( �i���ј��q��p>��/��aۻJACH�#BN��䀈�nA:��8��Bp���s��Y��E^^�.��T!�Y9Ar.�h�ż(hW�8x�k�:@%�2�&��2�up*�  �8=�A���{�O�
�k������h/d�E,�0�_ַ��(����|z$���J5&۠W����@�0P��=ѧbzx#���9j}ty�I˺��Į��w|�W �JW��N8�Yg�俙�v�#� ^Gі�D���Z�!��J���M�����⽵�h����������F,��?ns��XxG�F�������0z�}S]-�G3M�P赦�Έ�ŹQ�u�L��F�E��/���Nß	���]9Ĭ
?�4��.�Hse��J�c^kY������A-��g���
ya!k��U�YH��fh
5��j���t��o�D�B8��B|����=D�tZ��_�ϡhs�#��@�o�\�VNE�%�?�U z��u�)���,�p���s}l@w�����pI���CsKn[^��S��k�����i���V��4���;�����,t�<��M~�J)����|�(ɯ��;��_괋.�3�w�u�̚�5aggep$�L�:����#���jMB��]�����`V� �!;�@����h }��#8-���߬vW��"o��̳K*苊����q���L�[�Ok�HU��un�6�=<�Ɵ��D�Yt����Tql0>�{<rv�[�+(��ۄz��f�q~^�I��|�՛�&�`�L��O�i;fݖ#����\q<�H�4��'�K�>��(F�s ��<C�r�`�YV�>����)���nQ�.��v[ַ�Nm���J*�I8��y��ݬ�i!����H�5�NR�<����jW��u�O����H�j�L#�*cV@�5n��e� +�Oj���kUm��mx?��F�T�	��n%�PvM�K~s������ɖ�8 ��`���J���#��Kj�5~�f�Ч"�����C�P�<�����d��C]�	M� r�+�Ef�-��������g���3��aH�_&?l�@E
0� �ᡃk�a����l�a<�댦�<��7]?>9�^w��ҷ���.W���m�l�b�l�Ԧ(ޯ��iN7Ѷ�sۼ)�����{� �U7t��\�ԥ�2�`�P���,rÞH7��뛕�r������]��e�(���7�'��a�L���2�{��,-���U��1��88�b^��gʮ�������;K7˪^?"�,_�\���	g���@�'b���ql�KT�`@2�b^�]-b�t�xc���J5�h�wq�����y�g��{��?x���P���� �I�E�婲Q�8����wf��<�~�aw�1�8tQމ���u�7�*Oo�rF[�Qc1L��<ӻ�M�̑!���Nit� �L���5,�Տ�`�����=f�� Ub&�L�T4d��m[�i���s�=��DBPcӁg���9 \��Ddt�G<g�`xWXh��<*�GHE޾�"�ޤ/[&풂�I"k�x���-ǡ�8\Q�\wD\���� K��y'^�܄<G������N��P�#
t)$�H. �L�J�wg?QǄ�:�ά��+�d0�M�h�=8H�� �M�+���8'��y����Eխ'4Z{"1/w�����-����ff�|���-.��lP�`2+�+�l����˴~�~3l_OE�G��@���ח`��&;�-ZL_Q��i=�Oxk�����������{�?i8���G@�}�Z_1�vإ;u)��l�R���j[�,�^�+�����(H%:�;��Kq�A8{���YM�������~b��T���;�?3^�P.~�F��2�O�M6�zԫ
b˗TԀW#��e���cZ#���>m�E��~a�+n�?�Hܥ`c���-�3�1�y��H�����*d��
��(mہX2�cC>`H��ݟ��uzjm;�]�!�in��)iT����Y�8�ݪ�R�"kUKJ�_}�]��ǋ�;��(���4�1=��6>�b/��M/�PMs�+F4k~�4�m�$Bws7*���A����o�:���?�`3Ԑ{�-��'j������hM4���<�*������	�Aq2��j��Xo+�xT�p�_���6�ȟjVt�(e'�f��� ���P�U�z3��瀯hB`a�DSaӚ�I)A�kq ���i|���1������-@ɘ�@��%W�1��޾������#��%�_*�9-23M*^$�WVU���Gr�tf��vd���Z���u4�`�<u�gw�&�x2Oix))	(I��z`b�K�R���]�4�,�}4'�
̟262�|��q�֋o��R5H7�	�d�Dd�I~<}�U-;ʤ"H��w^��P�TP���>�urYЪZQ�%��Щ��u����&'�"����:�~L\t�~$�Y�?�]xSY�e��d��^�#WӴsQYw����m����gMq-/tU�S%!
���#u��|�?
��s��k)�1[��|u���ű�dJ�~Ƙ�����9��\�A��~{)�N.�5�:�4]�����H!:�F�\Q\,���?~�_1�;�t=E�̋֩A��&�mn��JqyӲ\
�perz�GQ)|kͤ8;A��8^�:�Ξ�xQ}�i�?,�`A�ǂ7�o�zz{R�rL@Bh��v��5��Tj`�3�A�Lt����bƶS*�]B�^�φ��4�*�7+X�(A��Y��/>�LҾ��������B5�L�ȟNά��q�.�C��{i0�fO��� ~=6=�>L����Ҩ{v��&�N��O��3�<;^�)�er����P�@������j�/���Ո����v*� y�'ͦ|�}�m��^�ͤ�F��J�h�?.�nA���d���e��-ʉ"���ȁ��ȅ��|�jՈz� ������}� �$�_�q�y�$p>�E�}��g;�$*�(�yiܰ�f��ms}]�ŕ�g�)i^3C9(�֘<���(1�m��]��gڨ	���.��%M e[�9m� $0D9[@�x<�	��K�X�j]�����>3�"�b��NXV���n:44��n-cEE�W�oC�z�2@�3y%���*���(K�nbw�G%T܍c���~���D��D	s����F�﷼��9�>���_wnyö�M��)�U��av���"�]�Q��=+ J�{�>����r� �p<�9����/�G��ۆ�Dn_A�����u�_�{x�^v���6���\�F��Df)�)�`�Πh%���]�z��L����R�A�h0�G�nU[�%��`C���q��?`ǀ.&e���oB52DOQ�cś��f��_jk��F��A�� �Y��ƨ�f5~�eH���~�Ɖ�\�ŷ����� ��*u�k{}	4K���zI�f�8yn��KK�Ow~�󎇡�O�F��E�y�/5���V� !��f��}��MRh4bA�D���ա�6N�2'vQR_���éÆ�J46i��7Q1�׭��j�Ť���y�&voxJ�:R?��ù )�X.	A��@����}8�!�{�`+�v,���=��u�V�E���b
u�E{������s��%%�K�Qf�b�
�����6~�Z-ӵ,��a��+N����R�V}�s2I�/�<X�*F+ԎR��v���;1P ��:�_�>-��D�ܹ������:�D�w�������wvE9��{�.�""g"���?��d��	��ڤ�����L%w��[�z+E���k|nr����K	��9�oGGޞ ��h�SmKv�Qs�V�6�
�"K�N�54P�!�S��H����0����7���ދ�h��tM�}  5& �U�<s� �zq���^��S��bO癤������f���f4�`5w� ��j����!�zR)UɱRY�#��=yHY� �Q[�Ҋ��� ���h���*�n�(e���s�e?ٷℚ��D��M��O�)/W���m}��+S��tS|fil'���	��*��z�J�9˲Ec�M�X8����vonة�(Ű�W"
X.�B�Sq�����Q�,cl/�-�{���B.�hZ��1e~�)����IG�����������U��s�ׅ��pՌF@�~/���:/�'zn̟���
.&�;��?��Ď��h�N���X��-QƔ���ř����Hl�F��6���Y@��,O��S��rh���[8�m�D3"�^�G�j�J	�jM�^ыz<C�^�(���ע��$)�rQ�gF������/K�j���*�]t�-�܉�N}�RSP��$t���1p3"b|3Ĉe<R(7=�ڹ�����VͼѼ븳Y�I0���<ǲn7���<��|�U$E�"���u��<[t���b!D(�T.{���S���b��4���B �$� sR���z!+n�9U�Q-�ڛd��G7���\,�X�X��kA� Zo��*$�w;s�=%^!�����=�f6�Ͱ�[����S y)�yQފx����F�gX��e��7���+uHzD<�Ƈ2������uX]Ce�U���lk���jQ�gI�%f�/t����ȱj�%Ѻ�<�k>Ji���}�����b\RK���9�U�-�<����X�2�f=m�ޣ|��s:�P����0_���V�R+_/��@?D��D�E��XPjlE#<�M�ik��Z�K塏hs&r�SEK1@�z�Ť*�2fPk�ݾ�������%G�aN�MW���.��m{�!�r�E0�ob��a��U�ş�����ZV�N����^g=��Nj�	$d4��l�05�uc����È�N��7T˦1�`R��{1�)ؔ���f�����������s@ϻk�ypn%��A�+��GKI Rt�a�����<4W�F���Y���/!�&��wgnd�ChB�f�/�}�&3Ʀ����#����A���b[O?��K�פ$���Ē�Ƌ��$נ�W��13ٔ١�&����ia^� gBxZ��Z܈�Z�knk�H��'Vs-֙c}.N^��G��W�<B*`���g�%~+�>�5�اY�}KG���7�q��J�I2��ȍ����m ?��{l4�\���t�v��R���E��E����mu��V�ug�g�P2��i�]P.[��+j����� :U�/1��.m懑����\H�hX�E~x�g��+���խFu:�t�
�84�
0�~e8�w
����(0�Q���[�/b�B�Q��
��y��^Tբ��~XL��ǁŘ��B����^��/�㻑5��}��d�r_�d���K���9�qW�
j��a�����#%��R΢�=~=�7��\{����ߒ��z�M�to���фM��,;Nn�ͺ��~L���KUfC��6�G�9h�ffN�r�Q�hq��H2��MU�1�b�B2t���Y#_���J��0#��[!c��3rG�GCj��G����K��۲Te��&؅"b��Py�����J}���ٻ������D�H���_⤍��g�.�fmO��_?o�^�M|��J�D�3#�|Y��3���p��1��B\J��F�6�d���4ΰ@����O�Qn  A����ZԽ�h���BD?�w����%+�D�&X<��*G�9�
n 	(�`���|'Fe{7��퉥=�՝��i�*�S+'#%�-�J�c���tx��viN9�����g2�������ƃ���\���ǫ�Ɏ�_�>VK>�멌���@�?T�<�.��W�au0�[�~>��#�%gg_�z�~�A��(l��ESg|��Z��{n3Y,O�i�vɪ��؞�0B�I3�@w��^�Wٹ�·xL?��Ex�R�r��d�� �&s�}��*�X�7�d�����i���޸j$�﬑�nTW��6�K� e�}��P}SC�g�D����R1&�D�� $�&�S&�-!�k�*b�;�@�g�m�Kc�gY�7@�P��Z��0KN�T��!�U�ȼ��a�̆�c�����<O�6���u�y��k��0�{�y;ר�ߑ�oak1�J_�G����C�|U�P�ه�.�q��ɲ��,�&�I�m\f�䧟�D㈡��Ϧ�;�V��'�%=��يJ���	<��)NV�N��ĥ77��]}ĪPQ-tA����4��N��!!9��P�_}ܕ�v�r�>=��?���ȹ��_7��?:���ny�Xr�6^��Ղ�X�I���@����^�˜�S�m�h����b��|�5p㎭�m���|�|���v�Ʋ�f������i�"�L .��W�g(���@"16��WPh �]Y����?:@G�½�6���^����B� �����h��P���Pڴ����G
J�������6$_s��bTq��/]�'��},J����k�F��XpX��o1O��ז����t؀Ѡ،����
���M�R'v5�$�Bj��֢�Z��"���cA���4ͩ0Y��\l�\����ߖ׷#׾�jz����Hj��@p����'�ǜ�ߘ�E�r�4��Jz2v�LV!D����h�>�I\b�U!U7~�0嚓,�3���!?��]39x�#!L�]A�ٺ%W]���q��!BX4S'�2Fn���`m�� ���U�� a3b�0�J�����iw���ǅ�}�;ƽԥ����Q'���F>�I�f�"Y\�Z�$����5f�Y��n����_�C�l3ԍp\�Ý
S��)�����4m}����#�`�/�T���pMd"�q��а1<5��ZѬ�a4@8cj���l��!@��o�,q�x�mp�mEGx�m��('����M���/��c���P�$H ��������ô�,H�ڿ�tt���d�CK����6�`�1t�"Ca�Vy� �-
л%�9����\��i �wƷߵ�I��kb[��N�oz�b�T�6����XN���zf���!�W}��`o6`����Z��S��y��_o]0���e2N���Պ��o�z����Xi֜r����ȏ�2D�<a��׺�^�����-xt�i��-��܌�΍ap1U��
�6وIb�F�!P��'S�kM��i�Rn,���!���[�3�0h���dw�t��>�&*u�&��N�������z��iy�@�N8�����KJ@	`��!�;:���S��[�[+���)��!O�/���"�����Gpp7窩�P�wE}�>�g��Ig����o��Mt�Pz����1�� ���+�}'�m�@��K��I߀^>��3�p�C3�٩�Aұޚ�-�	���$�QN�=���~��5x�����?(K�E����*`����[[\+F.�k�n�Σ��x�ن��ɠԯ`��xU%%N��?o���"*)���Y�`Srt)���lz�M���(�(���6�-؀���������
Q����D������z,t�4�"?�8ӄ~��yr�7�J��G��é���5Cx��0ϰ�az�����B�*�.>�(Ym��p����pk��@��( �d"(�s�M�5�:��A�z�p�j�wRǖ���;{������&|��NBͦ+����W�aޛ�r\ �=@tǩ�O:.�ӷ��ڈ�൳��q`Kru��PR�%o"�Ca�a��d��@j҅ir�r�ߩ��D�(@A�
,?�II��ϸ�\�$��T���.�}�`]����*`(��b)�؏������x2� �� ��:�#o���}/fp5�%!}�e@�k�{|��u�.���]�}�/�E^������	+���5�]���{Iw9�q�M�qֽ�A��1�=��y4���J���-�U��/�)�mO��YWlx�:\~n�e�4���Ώ��V�4�����3` ߰B��\C8ܯޚ�a��agC9b���m���A�H�g��/�+#�z��+�(O;Ł��@ՠ����A��J�͹�rnz��DjdL/t�{·H� C,8�[)�rv��/�9H�ُ��aQ�^�Nm�!휣#-�t�㬚KL�����y��
=�$�)�������Z㫑��pR�CX�y��P�̿�+0#�c��V*5oe��m���Fx�6�v?��+? �҈�n5�Pv���c?g�8zۉ0�F���?��5b�-'#�q_UTp=n�	BJ*��^&9+���Ua�H�Q� s�=���f^�$-t�H�6�(.!Ś_
ai�XA����e.�}byK���H�;,�-x��i<���&~3�5CG�E��N�ܡ�hI�?�
��)�dw���uښ���hz2h�0��_���ę��܅�2e�H�j�)2i��~��h��m����o	#O����s�}0�T>aIp`'�@���r|��r)���PY����Qn�{#1�os�l�����q?�٤�
�m�X�"N�#Z�Ci	An��k�RN�^�q�zOZ��j���Ј���O���j��BX(�1���|*��0����}>HK✿���gX����c���(*��>p�sn�V�X���P�LO�g/�̐��x]���=�ca@
LNq���O���lPO�3��Ü�l�N�C|M�J�e�3{��B���q�K$ ���g��h������9]n�� ���*6'�LHϙ�sW�-XC�˻�T�GOx$)�M=)�ң$z_�%]=4����R�"�`{��,HU�B:Lr�2QS
@����С@#�{;;7�Fb�_8o-��%�� �Y��&�@/�[�HX�����D_�����%����L��'� ῔C�N\]�s��A���]O�W"�������T�Ǘ�Y��`)7q�&a[J��s�.�(�΋_O�Au��K�ȡ�m��vɰ��9�c�=�I�Ҩ�:��o���ojR`��Ky�O�K��:N_9�	F΍93���*�r�����ķ����-P} ��߬l��cO�]'��@���R�Y~͂h>��G��e�t�6������Ƹ*+�� �c�DRՊ��Su�71q<zn-�Ձ� � )����,�:4�����Y)-�@ԏR,�A��h���.��ܿℜl��"}n$��� �;��6�s͊kӆ��\!33����Q�Y�;wi
i-���ܖUru��A�q�
c��	ɒY��7���"��Ҝ���2���%���B�洐7L�c>�p�xMV+��`.��4�K����7�dn-��f��יi)g+�1�R�P�1l��z��Ք��`�4��`����֓l���J7�������9}YL�7NyK��B) ��!��ɝ�fW��O����Mf�_�t�ߘ�k&�kxEc6f��v�拝r���*طL�e�-�_yԁi�x v�n�
�3�@�	m�mX��X4f�T�*2��.��x "H K�=!��ۇF֞\3/=��s�iBe�[��&
 �����9k<G�I	�/Q�8���Bԥ3 �e�vk�qwa�d�vM�/0yp@��]��1�C� -��ał=�cR����2��Mw26����Ҭۚ}��m�Ё���v8�XH;���wƢU��.摗>�y�-�7#��0�k�f�f�L�H�޿�w*C-��qg_��t�x7���C+�{�������H���P��{�ëB[�M)8���-p�4��C6ӡyz����JJ�`����x���O�y��H�(+�<h���ی<�o�~�k�[�,��1���[��(�z1u�tr�Ӽ��e���V�:��Ð:����hQ�q좒_�6����}�G�	�ma���1=2@j�����Q`��zD<&�CF�8CN[�#0��a�K<ߑ���=��'�;�O��Y�K���M�t �����c}��ĲI�%5��ް����v�o�!�@te�h\Sm�$ ׍W�dw.���o&��;�������>��9>�}������� �*>3u�4@�5J?ߔ���ϲV�j	*�:�YI��
JE�o�w�|(�G>d����]7�.��CYj�`�o��h�P�vg�	���]��[氡��~[m����vG�?L�}n�2_n�v�fxM&�ZC̯��ۉ����P�a*�\I�@�H<��rT�ky�#F������9���.��c�-a$�����1��ܢ�Ǭ ���J���;���|���Τ/�~i�('gSu�̀a:`-~ec ��;�����x�ѽ��Ǝ�+��>xǯ���'��Uk�b�2�G�ʺ�&���J���oO��{�bX� CV�,����m��t���iʧ���Ik��(�����a�hT�0���j���󭟡����/*0!l��<QF���'[s����t�B�����A#����6��J�&5X�'R *�G�̠�������J���ηJ�K&�ڔ+��w�3��6�~���+�|��~����A��N���Q(I�+�����>n1Pv�;<H�r]ْ̍"�����h��m[�R2_����b8B^
�$1`9���DU�V�b�-��
�7jU�<���>���?���MN��g�SE��'͕/����Gs-$	 ���X���^gb�a�?U72�Y���
DIЯL��#�/��#�O�Puف��6�¨4���]��A�]�KmEL%2���-�װp9pץ/��P��I[|'�N���ұ�������B��c��!��tM�b�m�I��\��a*60�Kb��Gci=�0�u��2�.w,t�~�"Am�B�j�z�!�;�Q%W���#� �m�d���p��P��u�Ql"//���t�P�;�5�(��|4���i��3��p��%��Ëh|�:�o�/������W�Ï��Si)����c�Є��Z�m8"4�r��s=�B�pЦ%h�b���,J��t}���~���ڏgY�>F���M�b�k}��uW�W���8�\�5�᭰�ىxm�˻&��k!B�LV�Q&ƙ���YO~y� ����	R����.��gV����ⶮ�w�Em8�MGɇxBA�q&�J۞�/3?����C�LF��cA�7G�<Z��ԫj���4a�сuq��<
��|�C}����Ǳ���}�d1p�vEn�#TI�J�R	��4/BZ>h�nf�'���f��ݰ�5;�7& (�E[��i�֤# ,�e"�� ��ï�/M�����s��y�s�%��g�A�m/�|V��O�
G>�W���YTn@v�\�\�99G9�S-� x`{�R9*.�\��]�l�e�%��l�K�Wk#�lrƷB��b�������?�v��	��5e�����4��'O���Hʝ;z�2g�.͛�w-T��k���P��]@,":�q�!֨��B�}�fl:*$U��|y�c�0;�!�2������1���9�ȱv��71��(͐�i�K�"ƃU�t4��y�	]��'ӽq��[�4���9t
���O̺��D�	N?"��y%�y"��d)_�H�P70%�j�Gf����Va����<%��|�P������0D�mp;���L�|ݕ�����C8f�tѮ�J��k�pԘ/QO$ ����f��臹jӧ�Z��:Ac�xӠ�A�j.D�5��%��0_	������%pKHZ~�r�����I��D���8�0"��l�X��c��X���}$�9���G���x��O���zo!N��Mq�.�a�>>Un�鬃#ji�*��j�PV��5�튋S��8�S�������`�8B����<(0v~kK����p��sX��A���M�ϳԷ���9�:�i=X���΀���\K�i<ֺ�>�J�cT��F�W��E�g��`�Р�/t�ѹiD���}�zG�+"�W����t��<��h�)���۱}6C%*��<����������QuPk�k����䙤��J���z�޲̭q��$�p��MpԞ���($̦l�!�� �*I�M*V��,�q"�I�'�q,��9P�X�E+
�+�*ܟ\�H���w��<O.}AʞE�C����E֖��\���$�}��˚	��mb��2�� �V��%��}�p��3�f�2s-� 	����v-�)���D8&K��6ke�JCd&=�&��ܼ�Ԏa'`��ě
���L�%QF"�@;`�w��ҭ���f�Ln.���x�D��x~�X��ߗl�������(����8�`A>�fD��ԡ��5��FX�}��2�����wa�
�9W��7��J���n�yǒHZ�6t�BV^�\�+ԕu��~1�Cj�3�&��
2]6���~[Ӕ�"749J[邱`��'���
)��ͨ�Bs"����4�X�(��޶��F�IeT��#۪a�����e	u�̡���+�/@�`f������R��7>�uH��4>U� |j��$4���\����W���o$�{�%z�N�Y���W鸰��_{�K�7���rA���}��ef&ȡ�4ϭ�cTG-����?c^<Ƨ��^�
+}`G`�$J�� ���
$b�> @��KG1%�����.�o�Gѧ��O�t���Tc�������3cM��N��[��LziR������4��l�(x����p y�a}<�.]��5T�B)7��ܨw�,�O9��R��E�=�D�^�1�u���兘K���/���0������Ɉr�笁��GY��UX�]NQ7>w���n�7�+�5q���_�F�9za��z��g�I��������}��Ѹ^36ؓ�JE.��m��(�3�>͆�	_��."+pV�@�.ִ�����%xz.���4�TZ�)ь�5�O�Ȗ����u����J��<9�h0�����Ah�B�+����0��rR���e��C�pd߉���L�)@�
Z�H���(o�����8�cx-T��b�/�zܰܺ=���v���"��h2�ao��"��^�W�e�f�r�v��V c�w�5��y_��wm�[��ط�jK|�Q�B��4��VsM�p�n�Ns��ګ�F3�ZE�i�r��:_���]�O�xP'E�a��25^���l+Q��#٦E�G��� 㶧Z��y�Ɍ�����et�n��+j�UZJ.w7"B	k��s}y5���ޱS�*b��mr�+d��!����f�h't����e�	[�U�����¥C8m`lpJ�~���<q|�{ʶlΞ}�by}H��.�oq�tII�oX�z�TE	!��:����A9��(!�L�)?@��wͬ��t�d"@��ݪo�ؿ����"5>+ɩ	08�ji��-�g�Ŗ[�e%c.�n�����iz�q���+�"�@�)��*��;�s9VK�I�9JE��5��Mb��і
DS�WX��[���7��O����vՍ��fJ�$��e@�r�Ǜ�[��χ! b��E��hP�\�eD׾�qS5 I�K�x�{�Ѓ�=�\}R[!.��}�C�{�FR�-�����h)�=r��la4[�	�Cpޠ��)�w �B���c�g�o�,:�m�Mⵉq%o"A��J9Hb��"+S���։!�ݦ��y���*����@(�Z�J�����?�񲍀�N�e�EB�?��<(r�l��x	���kXY�2��e�zg	8��J��|����'�(f�r���,DJ�2�����h�>�6݇��?﮹��u6^��F�~�Ev�c���4z��Σ��3���:8xl��M��r>ZO <1Fi�SnF�Kn� �������i����xL�]1Dɞ:$]��i� ]G���1�o�ݴ��6=�����#c�M@����TQ�6bIcJ�u�{����z���R�!`��IfnqW0h9쥮;A2�u���X���r]J��W�Mю�P��L�x�bV��7��
�f'5�H�m� ��m�Yjϱ�5����L���L(��O!����?��H����t���5p��qUta�����ƦWK���-~�5��I{�;6��bX�&�^��L�$	��+(g&7Q`� �P�r���Q�U���p#s8֍�!�R{z�����$P�˺#m[!�2�T#�=DEANG��0`9f璵���y��XzZ�834,��_H�*h揍lL�w�Q��o��6.Rҝ7t�F�a�9�:�����qہ���W�r��Ϊ������b���]�qA���q����RNZ��D�b�rʜ��p/��ӫ�4J�~���8�-�q���hF�wF���ޞ�5��e�_F�{���d���q��s0�R�}�$���/�5UR�f��"��T2�0τ{�+�]�?  =���uP0� ��n�?
d�=�ފK�o���u�4"���@�/�L�2t�5�9���P��-C��DA���	��?Ȇ#��p�Q��I�ݔ�Կ�ժ���v�:h�����a��N-����9Q:�
���� �[��L�A+�+�1 ��f�d��֪�h��@�B�-?Ma�����;��S��m0����ICg*��̥b��Ó�M�J��a��|��4���f���;%;������8�t�$�(l�/X`	S�ktJ�����_&�*��{�G ��D�^׀
��6����4"�W�ښ��F}�����eF����O2���C������H\|�L|�N��h�p�������J���^��4n�A/h�A�N*��S��B|1������;���U����E=#Z�>Cu0�SF�-m�.��a4N5�"�J~dܢS��_n�;Cp�M����^�	�<c�&�Ѯd��L��I�H��R�NR���Z �i;��zf��,x0��a��c''�[�))�TL�\[�:����B�aG_�B(5xm��y|��!��sv�A�a�8���ןI(\!N�T���Ih#l��6�����8u��i����� �!}�%<ï2D1�M��w�|Wa>u} >�dpA|�G��A�k�2s�>�5M��O�t��/��8�Y��ب���>�y���0����e�^�����je�0��l+�qe%�b���h��N<��ݡac�����[�sUF�ϕK䍢s���Ń%�UÐ�0�T߷��⃗��$<T�aAb�H=�@��F�6q1��D��_��@5.��E�ǩ^M�f��6����	˥e���z�3�=��p06w��D�4���(���,��^S������3�� �8�	*��4A����S����@�L�J��Ѧ��i�[:�t��������V�rmb��h���W��Ϋ������X�<5�W�$&��\��)c�Nnq�2�d��8;�X�}q��P�,�X�{\���d	�MTƙ�V���H���J����<("O���,��Xز�EnA����lq����[��PUX���N�*� {�Y��R��q�	F��~�[#4G)���!��"��{8ֺWW�� �,rYoj���!�ES&�4�I�Ko�Nt�Q��t��[��:��C�4VQ�$�l[���m�������-�tDn�ߝu����S�H��$q�~?�o���Ntp�$��VXD�%NWu�}9_Q6 Xu�\mK�ͯ��z�J�"=���l;K�[�=��{-�%\~6���#�����R1��)����ۖ��'���c��n�����" p�ֶD'�nğ���9o�s�\� �cေa�]lc�v]؂��ڰ]E� O��kU���� H=jG{y@���~�:?��uh��PJ�[Kޯ��0��#��X�����������M�;H(l�zE��t*��A�a+l ��$a-i]��W��
��
� bՇb儶m�ɴ�]Q��7z5���J�z��Nn<�s7giۀ�覻�AQD�*!>3��K�tW���L_o��`������"5����4dAO{��f=��6Gݮ�٪���z�Nq�S��nT7����t]�F^Y�����#R;�Y�03o��Ɓ�/K����^��|q��s�yҵ�"��,^0Rʅ�7~���z`pQkX�p �ʸ���l�d�����fE��#D�$��asu����������hZ�,����kб��,L�Nu�-� vEy�n���yc��GD������A�ݎ*��"�ҝD�=�g��_}�� ��P�z'�ʽ���:
m�So=��y�C�_%@́���cD����TOl�Vg�^�����6�Q3�T*}mUFǩyT7�s���
�DLەY�6$bE8�+��0u�]���	ڳ�<R�cKE&�9&ɤ$�f��*���Z� ���ԙ����J���c��&�I��qJ���x��XP��fW��u}`�K��^���!�[��1o�0�>M�;��TZ�_���� =<�6M���ϖ�����n���tW�=�ƞzx��k�2�\A2�R�I�6��*�E�U0H�׉�x��z����6���dػ��
� B/V��(�X��aiC9�����H_hu*������ѮL)�JS��#�5�!�,M�DK��т��+}|}�je� ��DEC�@�����)�� �>���.�����J�̕l9�49��%��E�*��_r."{	B��l�B*�ּڅ%�.��>Z�� ֲ`�����Nt<~�*���;a'�g���S�ny����:?�U�-c�^2���,�\��?`��(�s�V��	��}�N���������򵱼�N}Z/�q��Ujx{F.u�oG�-��1ս;�J�n6q7�14�H��^'ʂUnD�WW%�A�,�e=���6�L���`8jBI�b`ȋ29�-�VA���Մ=&r����]�W�}�OZ>�tood�T���m�6X��}1T��@ۼ~�)NnIo=�qG�K`�iL�Rma���R_b+�?�t��s�_'
�S>����,,\L�h��-�����}+��P%K;A��/�C��S��,k��6��(<�LB����|��H�F��g�%��P�s����o��z�澄$	P�zm���1���H2E�Z�Xr���n	���	�	ݥ*S�~��`%��$o�;W	�'��Q�'�1��gS+s`����ΓvUJ#8����z�ɟ�9�X�J�n��_�~�׼%K#x���NK[&#4t_��ڒ��i�.}�~�
7�����`��$h5��]�S!fm��1���]�0$��P&�&�1!�R��k���J=��Dr�K���{i.�nI(�;�1$CטwQ_��jaB�	�)	�a{ P��DU��K0'�˕���+��=s�L�o|�����e�(�n�ITÎC�	<n�r�ܬpX�ڵV+���G$w�ㆳ�0u��w���Bn�w���½����X��N%�Ye@�ck������O��� �_BI���<���<�UP�)i� 2��e�
���֔�U��1�pt����83�M"T�@�j[������!���j?��ep��X0F�����=�ʷ�y�+ą���TP,���:��x�[GţJ�!򥵵* l��˾4_{P^����!^a�
SS�R�ުV�.2H��q6q�.4�T�֞W��H�~;D��~�o̝��Z��F��`{�99֊`�K�n"��ݞ��:��W�G&,j�hG�w; ��DT�p��Ȟ`ؿ6��8���H9\[d�������U�"K��\���
0�c��I��yͅ�	� +�R.�']�e���3��������D�玹g�ꪪ�_�U����Wω�����ڧ���zG)�fݓ�K�	�I^�AX�(� ����f��y>3L��νٸ�ZW)?e�f]l3l^��yƆ���m��To�|�$�]1�"���l�ҕNRG��Y&_����wYv)���l;R�)�ۅ�q��da���M<���e	�Zҋ�p����7v�����w��ŋ��{��^�.7Z>��Kbl�������%Xm�:Z\��\!��I�l���>��7��
�,X�VN�Wm�n��>�;�:;"2<JN��n�H�X������ &���-!�m���O*r�ď������x�:���K�L�ĉԍS�/� �|)@`�5#h����)mޫ�R	y��	W�Y�H)��َV��%� ����]װ�Ӿ������
���_x?�ݥ��T�=]M�W❯��A���)��镍9Z���%��x�J�w��U��a7�I�+�>���?�+���M����]���Ϊ��pfY�|hUΊ�E���"������`j!���v5.]<���FN�UL������<:Q�I6c��3�e��b�UQ�����0��.x��1�>i��1� `�6���%m�䀮䥦�0��}0�Br�S㭘�,��t��>���d��[�A?�Dt�G�A�5B�$�4���oa���9���<��wt79���'5HC��O b=<��F}#34�0^Ѭ|.m�����`�q�:O��}'�3x��4�h%��lr����Ag�\pF�l5��hf��d*�
͖0#�����ȃ�Gx}�o`��=��&������ �#�T)�9���Ĭo:�Q��Q��9+1\������OEn�Om�Q׹=>mR�R��3���O6�-��+kk�t0���E�T*�rnv͌E�þ��&��t��Uco�/-���.�����n�{�OB�Ҭߋv�����~2�q��R5������X����A�(wLQ���i�+����D/~�n}����}�ל\!�͵*_���U$!%����^3I�4�U�q����;��&ҫP_���Zq�����Re�m�m���П-��P7>KؾKW$��ƴ�/z�݅����`�O�D��ܴ�.ڽ^$+�G�t=̐b��Ҡ�A�P+-S�e����'Xdv�wŝdg��y��>�1��!��g�M�m�&F�l�X�<7m~���Y�����S|��3�Тe�q��BD�6�M�T�|����I�u�KŅ�
�_�'�����3u�ؖ�D���U\��9���4��xXf�cˋ��6 (��?Qs��4�Q=�W�ܙ+���s����)��z��Ϭ��i��L<4�V��z��B
:� c���0��<_y),[
�[bQg�"}'�gXR��y6s9�M�F
��5)����Su25�U�DA1Qre�E�Q����&0�`��8��+1SBZ�Z
�ݠ�U5�)�w��Ӥ����(Ǥ ���v�����wa:�Eݤ�1�4dj7��!��,������%�rl�l5z�f_�@=�ă�<m�(OL�>��f���g�v� ��*yz�'�E��
��14�h��;�&d��>ޔ�WI$q�2#��V�f$���kk� q��"> 2vξzpںΊ�ƾ}pT�-Ă�\��a����S�����U�Ezo��2;E2{\,�}��W<����z�_��.v�l�[�E%��~�vT
���<�8*x��\����;"�nj߇��TT޿爦Ѱ� SK��I6+S�M��?J�a���
�J�_o����� ͵�.���4�˷���J�Uz����U<����пi�UA�9�^�3?�.?����J�CyB�u�p<V;�����q>b&Z ��?�j���2Q��(�2�W�}��h�<�	�/m�D��z;P��p��l��ݍ�ȉ�	8Wa�:yó���,��oFXsL�f}E��*K،壚;ҭ,PNI��%�YG�U���F����s�K�ؿ6��#@�	��JQ|¿���������U	%��"�{�Va�����@|�i�{r�oJ��s@����P��Z��a�T�����@fUau�x��`_o��#X�`��"�H��sG�Y�^p��-�qrԃ
nB�X
W�m�����_c�����Y���)�t#�f�#~�m��t�����yK�dhZxe#(Mu;(m��ɻ�Z�ɱ2IL^�`m���{c��1]bLxB�!:�lH*����[
o����S�#nt#4˝N��)*��B�����d�b5�
����XH%׮�M���ѯ"�Kne����+�wsiI쥰��&���1%:V6 \���q������T��T�Q^�B\�IC���w���{�8ع<�ŀ��Z�n��)�J��CϦ��~���s���l�	�k	���Q��^��T�:���[4�o��<����6�Ft�N'��C���g�b��@૭�_�̫^�'J^� 2,�ѽ�Kpa�P\^k��&M����|���r٨f��m4��Z�ިч��s���3�詖&�z[u#��ў�L��@6����2B�n#�� �ia�EV�J��#a�"�E���a&���)��%p�۴">9rx�ldC�G�?��L�܇:p���C
 8��� q��#��#	#�~Q�j�\_U��ǯ����A¹���`���KQN��"c�Em>K�_�:�'J��L���l�����e��+�4���n��Q櫕�P�]!Gmr-�寿0��J��gӨ�K���]A�r�]�����'�I^��Ie9$�|�%��?/�f�����V�����'v��#T���e�;��_��y3���L}�w�R�X7.{�C�+Z�\ܓ C�O�j�����ɑ!1�,	�QW���p*a�����|0���]��,�ɬ|wr\D4N=�i>ƥ�t�ื7��/swi���z��b@�����B1�f���A�5\.�Yb���{��~�^�{�e�튠c�gCW
���*�)�)+��8R��*nU�+�@y���{ch�� ���5��r�=h�.�#���
��Z1�x�ex'�(�1��8��9K���ד�{|T��p��腵Y����P�#�D�{�ج�� ~@�\p �I��=.Q3aq�y9��5oit~a'�!�`꬯�ÕT�0�/��~P;oɸs�����Ь��ڿ~ꓹH=ճyfauL K/�~IfT�ųm0Y6���m�EDҭ��3V�)�����2�n`}���2su\�:9�C��Mg�Z=��?���Ӆ�iAx���@	��#��w�Sh�!�7��)��9���F��Ӏ���L�o�;��yPK�J@�^����iO۽����� E.9�	�����U?�G��.��<��M�a�	������w��o-�v��ILӪ)�^�u0[#��A��a^� ˈ��,�����[*o�\p`�#�����r�:mvv�MΝR������q��Wd4(i��t{���{�^hg ���D6�]'�U�V��)Ӣ�"��jM�_�z&V��W���w(��oѰZ}���*�ۭ�H�B�?!7���cJ�{���2Dh�i�����̕��,�Ĵ�H�tƙV`�m�P�
`4�n�q�k�t ����̊��2�}�ҍs��~,f��Ƀ��<��'�Y&�&~�]OG���kW�<�A��jbk/6�R��#��~9].���*ҝP��˛��O��p�%���~71�v���X���A��8�������k��t�E�'�j���h��;P:�cIQv�
����t�����T�6N���aX.��C�oab(O/�/���+�`1��*�w22g�>�e)���*���G�Ux+���:���샕�t�+��	L���~����GyED�~Gq�?��A��&��4d3Ҽ;@���,�Q�mu.r�>d�ܛ�#P� 
~�����er�kү�f�;��F�n|��г�w0Ns�M<�Du�L��w��|�I�[�I��咥�j}7$�ր�[���[����AW����t�G߽�*s��}�����9s�_�sk�\f��}L�5�ʣ-�6�g}���8��,p�%`���2`ļ�"�O�L��?I�!��҄J�y!*x����,�>_ah?���͘�g�]!�q8Z,����u{J����J	?������R�ѴS��XZ��I�\9����e���N�k�	����F�w~X�Gq&|9�.��ɠ��9$�?n>VU:����,�P�z{��/^��U�b��N��w�/!X̽縵�Ha�w�����]o���:3����4޳]���`^2��i�ӓ��Q�0B�Sj�����
�9�����*j|��/��t8�eH3���,�8�,Ai��n�_L�������^�>Ma$TZ�kcV�B�X�Aݲ�/�P���vy;�+���z�N��� Xi��O��$�D1i��w�?���aN��b���w�o������R��/���&�nR�,�&���@kp��GL�¼����6�<������^�����,�i�������=v�N� ϘOx���x�,���N�C��36�'ek���4��'79�}�LB��H�<�j��$�0�Ш�[V_�')Y��<+�o�%�y���:|OރUB����3�q%f����h(��Yg�2h�q�@�%���ģy�v�I�U���x̓b�(3?��v�tY�L����R��[���)0�+��wIEL�����������;�e�2n;Tx�|��b�c��0�b�e�aĺ�c�>6��w.�`4XkfĲǅ'c��o|@��q�nM����"H�|��UU����؀�^��y��8���.�R�`�h��W�
P��V b:܂��)�WL�#�'E^��[��ת'��%�w�� .{��F�rf���:^n&�qo��<
�@���]R��S�\΃v�+���ak#X�R*e�TY��݇�V�7
�㺛���O��rl:�(�4՘�d&"���OĬx����Ϋ�C0��vc�����<E����q�i!��rgb���v������ee��"��C�~��d���~^	��v)�E��c�)��\�}��
���.��D�-;~O"���{"�]ph�C�мD��o퉉�D1��N1}���Fy�-�"1��h�{�oz �RL�㷒~�>/�3ű���Xy�x��V�G՞D� ��v9�������a3>�$�|��T,������j �Y���xܭ,�tj�l\I3�?x9�p
�m�՚�T�ֶ*�Dx�M�UQWto���*�x���6E�B�zj�|s ���H2)�Ե�)2TYO6-�Q���g��[	�UM~D-*r"�^՞�ޑ�e������^b���$j�Q[	_/��H{j4��CL�)J!cv6h��������nY���9��Fщ>-T����I>z;I�7_x&n^���Bv咍�2T��)�Vf�:K��Ҿ4#�(�e)3���_!M:(I >&5��<}~�Qs5*���]
���y�5����V�Z{[��I�9.ˇ���.2�

�,��������=���]�&������[)��(������
�N9�+�����TEq�u����%���3���WS��>�vb���-����٭���r��~e���p4��D����B	��>�@.m��(�1�u��qx6e}�te_��>�^����d�܄�Am�ue�G���P�Q����a�8aI[L8����;Т��~ȆGóNS�s5cEx]>I�F��<��;��m��Bҗ�q7�?���gfp�mR!�_���������&}�v���o��k���vF=^������E��!�M�P�V��q�/��?3Gz䢴�S�>-�����D��E�D#���?^)z�q[���$Y�3i]�� ���41���_4F�&�8�����	CB�bU���6���Y�f򐚗c��nړ��~Ñ^c�N%�<���D��h�yX�TM���ƶKP�J1d�GH�����9?�+>���9��iT6����ȱ@��ja��ꏆ�.�f\Y���Z�_f2��R�'��qD:���,GU� �:�9�e�L�������6	�$0�]����^�V��������\ c�"J���H��~g���K��*GL�k����xf`��66��E�~}e���$�I�蚥W���(a:��wb�z�Q<`������_��`w'��v�/
�������Di��W���H�Q>\099���K����N#��*�䡶o�@�����:��&��{w��$���|]��+3���nٴ�Sqr^�Xn�[r3us�	2���,d�C�,�*m����۟��^ �y&}f[� !�b��IX�]����qFJp�7�:�G���=��F ����C'Yn�䩿n�Imh{@^��K�՝�-!��\�o�B�&�|�+'�l��^��1�˭���QA��#���k�c�':L$�)OĽԺ��ݹ �hϔ��8�f>6X Sh	��I��]�#@��|��`� �M�]��=����:��f@Qc�ꆅ�0[�� 9؞���]N�99+ o��¹�c�k�;����/ݐ�Qq���O�X*꒎�4��ڒFANJ̫X�EE_�.�����zjE����C�"ィ�"��ub�￤X�6GRMM�G��B��z��.���%�Ε��n.(�}dKͣ3�F��̡�j �P����m��D��@]J��[�nO ��+��o�ѪA�ˇ��^��gn�P�2�%^Q��z���:�,hE�޷Q&&���5�"���31��q�+�T�Ǭ����,�W ��}�YK%��
���O��D'��m=B��'��bF��V���		*���l>���8 �K�{vC����Dh�x�z�Ր\q�{W��̀�`�F��-� ���xJ�ev�/m��W�-T���~�,ߗm�l	>��a(J�07�!m2Q*[��Γ�;Nj��Scz�%
f+�G,��y9��9kg�;�+�������@���"_+��p�s{���&)P֝�0�V�֏�T_:{�<��dp�A-sq*d�S��Z/)W/\h�X�
�)PG�F��Z��2S�5����[�N�UQ��=��<r�m��f�cZr#�2� �	*`��.������'�ui`U�ӸB�����fI߈�`�l׫���avw�3��V�l�_��A�� ����&`�` �?����2�������MC��֭ ��Z{�p��奭m��%��.�$�������/����� 0i�^"�[�<�������F};��D:�ol�|�q����Gz� ����a$9\��$Ĵ�<4#�3�z�S�rG|*l%��( ��\Ŗcj���{hQk~\s������h$�ơK�mݾ�7�m�]���:>I��������KC�?B�(|���3�����uVH���Q;C��dX�]�}�es�TE�cw	�t�S���Ġj:e����>�*���h��	����C�]�b�+d��T��R$�I�*�t�w%�!��q�V��\c�aL=�����~
���̥oo_w�� _�H9<Y��[�q�l�;��bc<X7�} ���G�hh�ȵ��ћ�����e����O�#S����ZP����r���#�s��=���\o LD@q6k���ڜ�K-��ey�fp���s�Yl�s�NV�޷y����!lN��ʟQ��:D����+���֑ڳ@>+ŵSGG��;�Ėʻv-O0�."��{y�La�p�,L���ȖɳD�~��E��֮����?a�l�@2��r=a�f��"�%z�j��"�o����i�q�Ӱ't5��Y�p�
'�b$(�w���{7+�89o4�YX	?+�b4fD��=U85�Y�J>�Q�S��GO(������J�C��Ƒ76�.����ڝ���/Wθ+#m���Jw8�5�Ƃ]���,���qt�([A�� E~���^���t�*���w%�b6L Q̤4�c��`B��tJ�G��>��q�z�~~�"�$t�	��nw���E�����%��-A-���2����	�)���=��Bܞ��8=� �2�;�ӯ]�/=��g�e�[�z��ȃZw�W��%�Zp� ���F��۵Q�8�%���j%��
�+��xk��ar{�����ce:�	%w0���&��+��2uLf7%:s�ձ-2.��jh����[�.
�g���e��[��v}��s�=�'� nVzNs�r�DtRZ�J�	|��Pְy��wJ#�/�3m�C�����B��wQS���:��K�
W�_�!;�h�$��G��[\�E�$�3{T���4Y���-��� j���9�@
�"-���a%ȍa��x������+>TkQF{J}U=؃~����9JF�]���n�3a:~\�p�3� bz�8,�V[�eG�W���q�Кcpc~d^�wp����di�	��i{ 5��A����V��$���#��S).���+ъ��{�4��`v��{��+����u��tw��%�o�ma�@_��+,�*K�m��ttU9�Ui��Sov��}#�'*�6:	��YjY���/"�d����	�Y��� ��/Aa���cX[��!��IR:ު�3?�w��x�����4'�4���Y��ƭ��5I�䉓�|V�A�������o6/�Fר��4\�����{ �n��V�i�Bb4�bY�8�kO��������LL�O]+摛���s�H���V��"|���0�H����v�Ꮷ�CJ!��L$��8��l�^�De�OO�`�g��8�A��=b��N��F�
�/��W�p���fBJ�ݷ;[ 0݉Ex\�z�Q��]i0(�@�w�Y�y�^�o�F!�}9�G�������@�]��p{ip��v��6��>4�������l�K���7����7�K�O����?,?�j n/�T)��E�9��l@�:t�!ɝ@7英Ϲ�+y�9]1�A�B0��������
q�D"�����lo����M{UN:��[����]�)�C��YdV�o�̼���є:��&zë��<:��}r.�xhM����P�( ��(`�+�D��}���}_Q`��^���/ux7v�Y䗑M��^wFރ/O�3����;g��e�g��Ӻ�A#���TC���q�Zz ������d�;T���7��>���vI��.��S�ti����&t����b���5��~A���(�߸8�Ga������׶%���_9h�R���	S2�r�bP :א!��E<2�{��q?��S�I����&�ݢ��/��V�:�Did�ܡΤ��! ��E���]R�w���l�(����T��9$��Ae������$�ۮ��S�Ԇ�����W�?��jX��"2��w�0�~d��X�RӨB��-ճ~�8d�f��s	n�QO�jv��^�+���Q�7u&-e��i����M.���%���%��;7ZCI�e������\���Џ���9>,�������O�d�Y_��skv)�s�($�G�r=,�T^��N[�wU�+^��Fˁ~챕K�������= 8�b���ϗ�gɮB}t �R�S��0 P��mn6��Ϋ�=YW�R�>�����t�a���,"�y���e,�h��H�H�(�G$9$-�~�uL��}�L,P��~+�����|+�No��a�.��Cb	���Ä��ބ�;q��T �a�r���"B�,�-#�b��|����y�i�s塾��S����͂ ^R5'�ؽ|�*��N�<��pB�֝�~�US@؜�Ҁ�����K�@Q��9��_D��r�3 ��*ZHh��qȔ�p�#D7 ;
.�jX��L��%�n�\��j��rgZ��B��l���{��������j84���6P��tOKq)����7�aro1ш���۹�Z�j�;�s� N�V<#Mb{h��_A�|�BRkP���O�$0km+=�Y���Ԏ�������/���"N-p=L�8��������B��gٱ/nq��*O���R �e,�8���㺲���({��
��lE�(L�sVb5�̫� �DmW�O���u�Wg̃
�˯�tv��\��&�25�kcԘ@��0���2A|�吵��Q)�jY�����W�y����L�qhp���K��h[&����c%���Zm�j�d���n���c�UӃij��7W���F8��yKJfE�^��u��5c��m��6/� B��Q�GX��ɬnk7�DBH��O왦(��.J������
K���ܠ���/g���n$��˷5�S��'���iY 7�r6�~a֯���FL�Gvg����,��4؀�m��Q����=;p[r��8�RpO���)n�R�t w�7�V$p	��~�_[Y��v�|�9|�t��.�>��32c����L���v$�z�d��̽�����m|�GRs��ױ��_.<Â�� ��zd*s�~�8����е+�R	P|�vFsu��>k�4N�c�Sݓ�G+=���W�G�%BS���b�9�ۋ+:��\]�[3�CK,Mh�$���IB���l
�������Ѓ)zb7eE���r�=,����-���9%����+�n@��A�Z4���+�Rk�	�,�5�K�C#�,��y]+MR׬0d	5N��~��va��L�-�M�>.v�|zn)e�5*����mP>���]N���:L�O��2H�Ѧ��H�*�Jq>�Y��"�����UY
�����^W�&n�A�*�	�	ЇT��'�(( z]���m�y�N�1�)v0.Žmƾ��c4�4-�q4=[�;�գ"�h��MG�1��ˠ�Gd�x�՞3�\�CW'���G��A�[�� D�����V�Yxw���B�K����+�9Æ�Y[��8�./k���
fu��Q�#o����Z��ʬO�{2�Fl�Ӂ��F�â8LTT!�9�4_����BY/1��.&�|���R��ˁ�K�a�Fջm�9�@�¡'�W��/�����a{
{</K_[Y)��-k� U���2���{*��g���h^���j�n���b��B�N*�lI'*� ���G7*S�6�,��/�ۄ��w��?Wڔ"�Ҳ�d�����z��������=��j�
�MvD�3v'7";��$�]�]�Dw ��Ẏ)%�K�ud���Z�wa&�Y�En� \�땭1Fox]���|�y���Pt�c�ό���;��:;E.D��n�5�48�����"9q����C\�h3MB���c�,��OV0�=��P-K����Z���d�9p)�2���a�.�)�4� S�����G}����?V�:�^v�G�	��� r�%�d�.��m�M���
�O6��̍��2���>�@�\�;����q��[�;�W*����}8��Rsb̨JQB4�U��+#(��x�]�<��KÁm1NE�MM��t~̩Lǹ��ͤ!�5t��B��5Ha�y���0Y��� S	����j�6.�I�Z�Ԧ�E�ކ�U��;�G,��5��S�Q����%f��n��Z��#�A��~�N�M����&�*P��X�wi\�d�(����@&:�f������8(��C�w���-,�з�����38..L7�/F������w��{���	ۯro����Un�H�DQ(��;`�����X\�GIڨȋh23�t1���B�,�D[ ��\�`���
�HUqHB�Pb�W���R���#�6~�[����U���\]h'�
y��?s?/npŴj�~H?�>_ߠˏ��`ri��Y�E���_�d��e�3�b���Bd�=*�v��]�2��9�F�H�Aqi���pq�����O��qb�g�m�QU�3Ge��C�"�Dz("��k���I۽�)�w�w�`��Mn���\��V�iȦ0��G^|]���cP��RG��`���������\���>�"�@A�)�W�e��`.!�A_�����v���������ˆ�>5Q>��o�Yqt�����-�8��f�G�haP'Z��V����|ʓ��#�k9�%���v��:4(����T��>���PG2�5��c���2N6opqTD����<�%���1%�,�C�lr"pO��!�_w|C�
ʇ5�|0;���?���o&��E��'�{7e)jo��?A1w��Z�-�+o�{�!�Bw�G��Yxz��sIG��W�r��w5�ˈ��w�%o;�i��� r�S�\�ᶕ�b�yj+�,�^oaa�iaO����5�^�$�dK{*B%r+�wn�[�yk����6Cpw�g��B��4�vx��e�|4�����Cf��UX�Јٲx�ɀ�䞈;���<��%��8w���I�.`���m��"�-4]q�+1�ex�Mɚ��aU�Uσ)`�u��
��<4ܒ`)s����	������i=�R`��o��!�?��c��9+������_f�H�"~*!��x�f�Z�g�n�Vz�7�!|�A�#� �<�#�ײ(�z�<U��z�P�F���`u�>���x,3�&��2�4�z��Cg^ΚĊ�Y���?M����ֳ�c\V��V��qr�Ο��o����oE�R��V���AU�f"���ņa��l�T+����{h��$�c�O5�2���(u�I0l��O$��i�>gG����s��=ҊNA�V�$��-���#�SeRK�0�t崷����Ϸ��7��ͪ����r����p�N:�u��m�Y����w�G'��A.�X�Stc/kؔ|����\NK���`���Dw�6A_$�5+ЙV�	gW�o���}d�6I��>��W��.����j�O�8��x�>��f�(B{k4#/�;�Q��/�5�ڇ�מ�n�~8h"�j1�^�pM��Ȝ������|��H��1����9��#��_z1�$���L�r�E`(l�u>4-9?Nnpf�`��[�wAk�up�,DQt��ȝ��u������٣J��B|�D�ߢ�ف�1����o���\1��J8�	Oi��e�j���gl�x1�f��"�Q_ɋ�/"6Éz��N��Q�9n�0�j6��<�b��-Sjy��A���J�-� k�;EaG2�#p)V��(��/N� ��t�zIԃ�d�e�������y���?$w������Ƿq�e��5�$�σ�cƹ�}fUR�:���&)FX�̔�?�BJ�mw�ŋ(�c���o�0�N�d��H	{VV,{�`USw<u�7S7T����0���l�0���(�Yy{f�_a���芛8ʇ��6���iARg�al�e�W�,վr#Vύ����\+�r��¸?WPՔ�urѮ��X��Z<p\�$Z��Z@8 ����`���|.��9د
�]�zk���5x*��)(��ǝ�ȓa�_��v��لP}��ʡ�v=��|`����2]lݶTfS~l�P77§�(�o6�1�\��?��j�XܵD�O��+T���0�CRI���$+��q�j�A谰�~���ٽ��~�S���^�}w�U�� �z���.+]U'�$�ǆ,�H��2�<����ڭ+�4oX�p���������Q�� ���Р��E/q/f��W;�y�fث���H�7Pt-'�ڞXq�	-{��u�m
���"�-h�SL�y����>CC��GS�� >�S�VM捣E=��&d�7J�9V�@F��K�,�%Uؙ��M;�y��I�g\���[�6� �9
�d�.+_<���O�[&3� 	�dDЭ�,Xc��I�ýE�H�l��u���Ey$�N�v��ş�#��%P���ͻr�[a˓T�]A%�t�"e��n�6C�$/���ɺr��1�[�{��*?�I*z��@���0��F$T ��fȆ7��\FW��8gJ>=�4�El	^�z��BM;9rs1���Ư,&(���� ��ߔ8T�F��*�����ɔ��!�ҾM�;�2��~�\��+Y�r�tN�Z��X�_A\g�K8�	m	�m�m�F!�)1����{�}�\���˼n8�+(Wl�Ⱥt!�
z�#R�	8�P����I�M��r�����.������"�jA���IJ�'l�C�g.�����5���3�M�m�#��Q
�e���"�V���_�:��vm���L�k�B�\�f+���>˝���,��!�����9��./��8������G�VP�p��:�ы��&~lE����~�����q���{ Ug0�"E"��w?�.�I�PKG|�"6�E��l�K;HY�_qyl�]�-z!�y��'2T��yW���i�p����TY�[5�G�n��	�S(�6	6�������v�]-5�v��i�Ԯ�K����,w�8�k`k$�a��R�w���ĚT��xL��Q� �Yi���a����x����_E�yS�ck
M�v>Y��_��T��\Fw`��qL�.K\QA/�D:!���S=�e�[>O_$O�����<'~���V�A+#r��`b�n�(�]�i~w�B8k`��e�����aV��@��
t�H%��Cdh�$_�C��]��-�a̧\	����ǰҸF�����i����,UAO��bR����,&&O�^G��1�m�0v��~�q���$��0��ym�s��r���%�P�M
�T���3��W9+&j!�c�<E��t�"X�%�c�G0�q�B-�W:$F,�D��,�2��}�����
}����@)r�ո/v���l� ��I+	Z���]��|��h`��k΅pC��V9t�p�G0�<��q���ةg(B�-��;YѾҭ�ww�Smc[+�[	#�㢟���".�H�Ǭ$Teü�;�\˭��{Q�Jo�#��ط�+���-T=��n�KP>���k�ޭ-[H�!�l��?�_,�i9_&�����¹��e,d��ʃ�j�tz%��-��)�k�z#jO�ָ3<�T*�<Usj�M�o[O&��d�{�)J��G~g��dkG�����p(|Vd�K�Qm���
��+V]�=�Ar�QԶ�w]��e�����Y>��s�Z����������nc�h�}!�s`�˛����%{R��(9�R���T��z�e|�5�NZ��F�9��;xH�O�P�F�n���g���Mv�|�rh��^�����@���q�������HPr��d�����_�_'�Lg(}����q�mw\k�����}�\����v�#����9 騇i �ڍ}�������K���P�����'���/�tF����w���:.~Nk��~t�u�'��ʿ��C8,���(���!��ػfJ�mD?�i��V�zU;,�ژS�l�c�-�U��i"��at����q����s��ڍ�5�Ò�L+�%�z��°�[G*�}���M�S�iˬ�����f4�BθU6��fvX�P��Ϣ.~J�����Y��)��j��'4�P��b��[H~2̮��cȯ��HK�e��լ��q���ݠ��9�����ˈ�����7�%�oO�&a%yS;��8�$�x��l����?�R:[�L<{��k�1�`����U���ѨF����`M�-9'�/xM
Cw-��I��V"�]Y-��dۓU�L�S)US�������$�h���!\�RR���5�l�,6���дn�b���ʆ�gY>M�ѿV�����BJ�)�l(<��g%���+G���gЩȧu	�&U������F��Ti�����eF���ŮW�^lry�I^@��Pj�(ێP�݌4��U$��a����.�����d�+�%�!��cEݏ�KxA�d И	F�L�S-iud�&��ՂQx�؆�30Ҿ7������	:�>�F=�d�=<4�vS/յ2�����Oɳo;֎_�v�E!���u��su�Fx����dk��ϓ���gM����s/��	�]O�0��l��%�}���-��+��.a`A�a[�Fe��?/`@;�U���v��`7Be��Urjn�@��@��t��$(l�*��~l^հ��->�.Y!�>0�1�8I`mJ�G��Q��G�	�@�q�k@�f&��ł������j�:0soHA��~{=O���Zbɕ}��րp=�Zm^��U�>m�wD}��~�w�?�ֻ�׾���5���ZB�L���J0W�cih���5x�_;�w�I��۟ xp�;	�{ڏ
w0���F웬<����bC��]���b5��;�a�w��3��c��"N5����Q�#Lb#ӝ$��s�qs�n�*Q�X-M�G"!�J�V�Z����.!��jeE�j��)�%���9�wb�:F˵����MΚ�3
!�����YGD��\����LA��h�l���=��~�{��`x��Y��t«u�Wں�q�XiXL�9�N�>�˺p����Zk�����\W�u���R�-��\��Jґ�gT�o��*P.vy����Sp��6;zp_���aa<��� ���}2l����T�Aɇ����o�l����sIK&t�&dj��|m���춣��X���/
�i��^����B��9�#X�9����>��竗��\�g�
b��K�ޚ�nr�v��z��/�'�te���aH�)�df��w|�| Q�?¤kP���Fl�E�%�����9ȝ��;� wʱ_�9�{�E�P�J���ȟ��Y�$�D�q�%6$G�k����ngݟ�fz���e���+�����+�i�S&wPNb����t'g*��S��V���mJq��L�/�3��Xt`z��-�n�:�q֎�K��bs�m�q/.��{#�>�e�yCt�X	��a�����h�R#�W�*���6��1�~f`0�d��(�ʍ���PЪS�/4�}1fčLꥑ!��x�b^.մC�G�T=��un�p�0�#��GHG�'�Nτ���_#��|�ܭ :��`�*�^_ѱ#�^uM���rqg̒���]��s�!��br34���_{���y;Wݙ��b��X�2'~�G�}���#綱U���i�	�z��̆	\J��B���d���n�P�V���z�r�Kx�+��D�?tG,�!!��k#C���F��Kn�3���W�'��`��#�Ψ���UYf��Y�v�P:�S��yF"=}(�l?a�û'�|_�X�A���Ȗ;����/(�Ti��Q�Bg	�A7.�ä��;_,?���#j0���jfפ�	��[��K��	�v��@g�;�����R�,��SH��N{�c�6YWͼ:��jBԑE�ټ�:�ҏ�Y���tοfZLPQ��y��|��j�;cA�aCI��	�c���*]�A�D�ǫu�u�Q�ץaxH}�<��KXo.��=w�����E���Z6�|=%�]ϊ���m���|��Ґ�� ��E��O�"��f�W��Qܨp�yWCה>�r�o.@~��5�D|m0�*��Ԡr�*�� �J#���o	f���:y��-2lSu�1�^zIU��us�vL�1&�dxṇZ��˸j}���5ѬD��:9�cJ����B�O�fR�*�C�$!��+M�Q�\y��=��/���/����A+���xntVos�������kx6٫�#�3�D;�~TkRH���6��
t���[�"]&�l{�TxҌ���9'\<�h��p{�
�[Ő׽�LC�fA��E��
��Щ������\=�����S+�B_�t��L�A�R�7�-�VS�F�٤j���lF����c� �BTD���ɓ('fYzD����c���'s�-���U��7E!#� �)�`�Mr���n����}CDK���^�K��`Z���!�5H�����}�����"�n�^^:��a-Fa�Bp�~`q��'�@�� �G�M�����m~�T��K�_����-~�*ZI��]/�� ڢN� _�^ߐ��jon���!z��j_�,W:<L~T�:��ă�cCw7�T誱<�]��BI�ݐq�Je�PrTMݞڞ+���A���aR9�0RK��!��|�ﴪי�4��Rv������)�F�#�6jC�q��%:���@��[�v�,e�6c�g�y�����:@�(��b_@&H�V	�|rL<-<���N�-pG*)Zrm6�h:�j��Q�^G���o�l�%3nS��lB[-0�dT���y����#T���}��U{L3�:�&��f.�BLT� 7�rT��?ɿ)����Vl!m�;G3��e�z(k�=�����[��A!D� 7l�Z�:�'����$�pDR6%����[�@�3�c�������,.��|�/85,4&������ `�"w�<����~,iN����6'[E_/_�Áw.G�P3�G4'�zy�4g�|�oRT��?b!�	�������Ljc#�7�z�.]���8/�B�$����-�T` �Y�4S��"��? c������x]a`���CL�D�X������D ����atQ�v����|��������B3�z�h�2Ww���� �w�Q���+2�h��R�|�6�_5�'y1��n�ǇӔ��8��X<��[ݫ_�J��ǳ%���(��B/��qd] �O}Ló�Wͮ��� D�k^��S%�t��	�;@����q$��P���0�@�?���ȅ���Nbu��x����7zz#��!�_�Z<g�A�����A;[����;{BK�u2ۂ!�@��}7>FߤDt ����w��h�9����H���u�#�.op�!Ӷ��Nh*�K} H�|�\�M�0�^�zF4>�����Z�΢q�Ҧ"`�x���+�n�d����W���@*+Ȓ+���U��_.��1�ِ9���E8ן�u�a�z����p!����aU3NiB�k'����VI�ߺ��
D�)��X��v�%��y��]2����S���'��>�Sn��K��5�D�A[�m�����"Q�Q<˹�xۮ#K�X���M��>Cםy�F��s��h����6����ya���5�|������]�Fp�\W��U�ϧ�@�q*��E�MX��:锻���т���7��w�<�V�ܷ� �7e^ۖ}�nar��=�o��c�Į��Z M�����4�$��fe��È�r�/PY��,��?O�A�����=g.<km�TG���5���3�I��{@�Q�9�G�(٥?��?���	ہ�%����BYj*�'fEu~��?AN��A���#��`��V)M�'= ~/$K��b"(#U�<*��C��g��4�G�G�}	�B���7	`�?�I�^>����F���rȇf��T��.����\hR�15�r���S�-{46�^�f�j(u�_���:6ҿ�q|�jW�|	:�9�h��T��t�8B��cH��K�N��C�ϊ��s����s�s�t�jR�2�9	V�����R�cO�ߣ!��������ZK���T`흚�l��'��LP��R�m.j�Fo�����?�!1��(����FD��*F��6K��y��4{k��h,�����2W?�W�7$b�xl�Q!Ѻ�l5w%��H#��j������x��(@E�Ĝtf�ƌ�����Nk������r�?f���q��BGR����h��ΒLOgTW�u�F�"0!��!�$A��VQ��ݠ-x󵀷0�U�}��{�U�P7���i�)"+	Q�u:���}N���p@j�:�Ƅ�@��#�f�1�x��VqMkkt�~�N�g["�R����ɮU�/����U"ܸ0��*GT^>Xi�I1m�d���g.��hʆAS&�w�m���B�5�U"�|�����qY2w�P��f�����S�K�(���pdH�6�0J>ң��|�u/��ֆ��@��1��'����= ��-c��\��Qw���P�Ì:��d�7�F�C']�Isو�W�;X��u3K��lM�"h�h6����$4��-�Z�����YVF꓍� Y��xec��C�����o��{�]ף��^%H�Dd�9��s��6��BY�?'��a,'6P�����9��vf%R���+F�T���M����*16%FE9JO���W�Vl{���o���<�c�&�h��&B���p�[rd?�����_t��C���Kg�]5st=�L8�ɘ{S�
.�䃿;�7"N�`�:o3�-�\��XY,`�����?�f�h�ks 4�N}�^�]�ƄUy�C�DJ4�����ޢQ�� �"�qʼyl�C��f&̠W]�RQ�Ss�Vڄͧ�Wn�d�' C�)�4u!��\l����|��;��k�M�����L�&i��:W���ft�d��/���0O�ɝ�N��j$>����|�g*�&�����G
��"�]1Y�����
�=��v^iU�&mI���]E	����$O��f|N;���<X��Z�pRy��u�q���9[�2�W�{e�VWn�,�T)g;X��L�]��ث|\�([r���#�v12�$�)kω�������y4f���ic��iy����ɬ3��S�����UϢaGjT��EQJ6/��9+�1�"]�Ϸ�'s���?�N'���k�s��'��hW+�+��ѽow�h6��&뭹���R�O);�#��~y����D�=�1�v�
��Y^0�kmEpX�X/S�5�ig]K�fcM<�� &���kq;��5o����Z�w©_���R�F����,W6���0���>5��/�7�)c �R��g����Lx �C_�sS�ᴡ;8.Fd�6kAq[0S���\,�"L눴M(�F9"�w�~G1:ż�D�qO@���\�n}���K�Va��Y�M�'�s�K����6X�3����_�"no����?r��4>�Oizp�L�����y�tˢ=�mu�u�f��ʰ���=�Ċ�]�&�ؽkj��} ]���Ȟs������V�	&p^�{^� *|�b*��Ϋqlء��JGm��h�Ah@���neR��x~�mhAi�n�� ������(�@ 3�&��M��j�<���y�F�q3���8&�Y��f�$�/Ƥ�b����Ɨ}��31��pT�g�1!t${����U���t&q(a�=�+f����Z�.R����oq�BX9����OBK����:�
�}�H2�ݔ��PL�ؐo�x���dz�u�1���p:V�������t/)��-:�ey~�\�r7��5Yj%���p�'�oZ�(�D�xD�1�r*�	S�h�U�����9���]�����n:=RZEfu��)GT�M�z��������S�?	?��0����H�6��p�ن�����e9�Ma�>�R� ��yE�<o{�9V�'���lҋ��[xtX>�n�&,B����M��;#�
n��~��v9l,p�ZE�N�y\+�/��?Q�b�����ׅ�8�d�e�P���Z�B*��k�|�@=@p߈�,�wy���X������m��kق�-�!x};�%����&��.0���9�g�Hũ��U�7<��4���
ܢ��m̶�6Nt�2���f]�Qt��q3|�'�F�"�U\&��6���'��j�A�0Y�\K�91��!���< ��]�������Ep�F�~�0��ARK��G	0���.�V���nݩـS�X�&��Gy��
�~pu�^ʵ �/"��Ou!�SA
�J��3I��@ �\����M�|��T$��,��Kx�~�]�!��}�k�S�T�(�|P��m�"-M|�#b�6��'��.�H��ƶO�x3�^x8P�筲�ӓ"�_�d�9�#*�,��N��g�;�۾�= �	��SKY�Q����J�24@q��j�韒'��a��]�*l-mtE:Xj�(���`) 		=u��"�תU������_��T��l��_1� >��	���*��`Ɵ-ZJ����#OW�MY���/� D�s�r�Ve���}��Q�A-�ܥgc�T�6h�G���&u���/�Vx�n$��;��~��~q&��R�f-��%"M��ԝ����W���H%��� ��ގ�q�����AyjO&��ɓ�
�>L�I/jw���ú�y=7�R]��^3(�*�
���^�@�] 5e�c�+g��ud��o��������̙�F?�R/!�k�P =����#�Z��`d�K	֠�fɵ,���n�E(��	�PV!�ϐfX��A�L�c��浛N�㳥����y�3M��6��������~I������2�^�~��oIQ�{\?���F�3o����{���o�t�g�z�.�I4�/�����ULǀ�ct���>i����|ۑ�Vmj{���& \�Z�&u]i|"w3a���
����!,O��&���sE?��-;�gP��s��U�)M��|&W�~�T���B㡻�$�6)uYTZ�۳���z�h�Ro�PY�R�^���@A�p)��e5�~�ү>����ocY-���=��2�P.U�d�s9��,\S����|�y�r�Q�Њ�	i&,k΀;�r��2y�P�v*�+�Uv<Z-�!3�e��S@"뷚	���$��ώ5r�^AV��"��#���������pl܁�����a�4w�KP�z8ߙ���.�)�iL��4�H��}��qx�5[s%w���~
$[a����JtE����)��yZ���trÿ�=��9}���,�b��(�y�N�9c�۵�n���<u����_�[��r�)���>y���9����:1��9]l��7v��6��?--d1ɢ#��ϭ���dM@(HUw�C5I��z�5+S@�}�ӿ"g�3����U�B{�C��6��qH��iXS'sj�z��
����ݽ�Z��yg&�q%��e	ʰ��A�b�������J�n]�~~d�����|08z��GÞYI������U�'RI�H^T�����)U��ߐ��J���$����EN��n�>y�]��v�C�抽G:)��S��.�56�����P�Y�[�1n��P��Lfݓ� �	c��(�HV]����Q��D�&���\�'��}5��[�<��<����vy�7��<�
'��_J�9?�C���>�2vU��U��o�7@rVb�	斆�Ԧ��
��%�Jt�#KPH�${�z�X��/s��Kű�|/N��o V�J�Q��Y����q�C!޲�opd��o�$��'3��t��R�@J�he�X=asy���:u�(���1�7�,!?h�Sq ���4�k��!�����N2��@?���<�Qż/��d������i_�RE8ϼ[$�m���6���V��&�|��:��nK���Q�tjuQO�̅�#�4������V��$W,bp�����ëG �� J��W����W����3t^?�
H����B���sA.��\�~vf��,$��,9��T�yV�䧶5�@���Eߨ���
Fυ���}��24-% 烙[�٠�6~Z�~����`�OW\�?��,�J�0D�OUڹXR���$Eg�����5�<����?A@�J�]����+�ZW������.;b������(�|BT-�<�n��EF�>Ҷ��"�k����R!�i$+n��E=�Z3,���4���K��wA��&:��j�T`�e�3��*TX
�L�壸Q^!�8�e�Rغ��o���"-���v ؂�Cn���_�:w����m�r��1Sy��pj��<�a�<S�)#r��5d��7���록0��QI�Y������*M� Y���Rq�E�I�N+�vA+��1v<��8�E	�贂��ͫ0}Kw���|\Sk��;5a�JY����F����N[~�p�Ȏ��kG6�8j�"�K���!��J���ױ)��$ܮ�KA��yA�����>|�����}�1�v����@�Ĝ�o���!�a(X�kl���9�$��t~@HRS�=\lx��)�����>��o�f�z']�+�o��~�@$�I,^}-���Z+������։*]�n�ǒ��=~��6�ޓ:Df��G8ncg��+��뤷崬eeD��rIHSo�9u��	us�'ݐk��<I�)��TC�z(swo�{�P6Co�?]r���4㥚�����9J���o���TC�q�ZG�|�P%�ќx����G�`����2�_B���pf�!G9��A�b�6P��f+���sB�1u�솰#xQF��י@�k��2�$�%�N/q|T�?g��y�h���w\��c�	S�4��Bu$Ͼ�F�� �W�/�Վ[�<l�@}�Ѱ�4�	����� 㫽�Ǹ����K(�ڱ�P�6+|s/~�����KrOǐo��r��E/�}R�9���7Ѽ��TS�s+���.*ٕ�����IM��U� �li��U��`�ɰ��Q�e���b�\2�$���Wx�#׾dB��1�`��#��1��O՘7�P��,�����!�h��&3�w�}��f�wY�<� �����H���=^��Y���SQT܋�哰�&I�;�x�˙��{�IӤ'$�W�Р�O������j"�~�����Q5ÝqA �8���?�k�ԁ��}W&�Plg>��oS�լc�)�%1c�r%�V�Y;���COf��nRb	A"Wq慩{���"��)�u(��B���$7\�$���n��<5I�H�n�7�|��|��8�)�BC��y�\�_�Q"�G�$�U�zΑ��4����V'��+�C�!c@*�ey�/�pR�u2!]��R�����!�Z�K��:`�N�'`�}g{�Q��?aZ|1����q^G��EG������!�	?W�ս��63e�OF�ԑ#Pq��k�8(�H�߀`���c��;��W�R˼�x��Y3�P�?w&�  B��R0+@�� GEWӭ?H)+�m2d +�:p��J(��!xq���3�����ֈ�RPn�L�|T�s�i����z*��G#SY@�;��a��Z�$�k&�iud�>�{k������0pH����a�������Q��؉�u4}��[zX%��t�V����W��>��,Ӗ o��:�g��u����47��z	�v^-���/&�I�����K��A�ff|�d�;O!���ҦEW��T��uS�D��b���� �S�_!�*�oق�������?30Y��G�b��E�#��8��T���3:��d�Om}3[�d1���+^@���	�� 3]���AQ�ҿ��6��GIᐈ��_�h������6/w]�;G*���L�I=�9 �׳�_f� �V#��ߥ�>ɧ��!h{�^�]4���}q�;ћ�},=�T��/J����ṳXGzM������F~N�L3�H�X��%�y^�OU(2������y�7�����&���hN�EG!}��r��^cq�'�by#]b�����EHB�q�8��1���d#��)p.iN
 j||��}�(6J8Ò�0�ԙ1<�o������>5�rs>�t�&�$�xh�D��QXE���R�0b]�4�ß">0���a�1�*�/�h|"�%j��_UQ��c����x!D�o.f[�)Z׷	#H��q��/idD@5MJO���l���gJ�Y�!I}�6��� {_�{�:wN�Go)��W������ma�?]z����Y�^�%d���[؇��@�@�*�r5�h���.e	 �"�v�8~��"���k\)]F:&�:��� 	ʝ�il�B�zۗW���C
qA����F�����{�m��cR5���&�s�م�ԗ�9lI�9����)Z��ƒԧR7�0q��YZ�;��V+��9]����,���H��o	YBL��0�M�6��Q�)5�8'2��Dozo�<�ol�	����`����1-�k�Ǖ���6]��l]��A�q��(,	1+a���9��R�� T	7`q7�pQ?���i�Y?#�P��4�h� ),7�Iܔ���5�-'��5�-��M�����A߬��$ܣ1�adF�ԯCRN�w@aI��m����N�'HK�܌b�<.�0�4���'�[m��-��#y�n�SZ����K�]��C{��i�����&�!���ɳ��#�Ic�(7�U�LE��*�~���AҶ������ ��@�sU����p�_]0�+�ŗ�r�~��k=hQj�j�$jE��u
R܄ǟr�2��|�igt&X��j���jW�	�{�Y��;�����}`����4+K�޺U�5Hw��h�-?�n��VBU�*#�Flݮ�l���c����p����aIAIӭ��c�&����$��#�$�b�^���k����<r���o�^4�bOh�qk��n4(��v.��A/�j��8�;�^�e��z����,��P�u��c{�6{0�A���D�ݪ�\h/����+��2[g!}},�?�_ƁN�L��0����-��wmu����Q�e�ikL���W��"���q�i�`�6Y������<��Kk��^������`�5���q%�U%��	�����0�^�9&��.b�&�N�@91[��������w���~��N�*�=�K8�UU�y�V����vx�"%�[���>E1�	��y���	�v�YxX��\�:>es�F�G�6)!7Ȭ�0i��	���o>?���s(��j`J����a`�뢱�#q��4��bW���ɾ�"ߘ���lj�u`=�j�8�3��/6}���c�u�y�n]��?d�d":1n~��H��xH/�G��p,���w��GA�>R�s��wV��s�W�tf��4�H�8M>Ћ�wH�ovۓ���B���9�*G𥩧��&(.G�)Z���E?�j>0GU��o_y���e�Z�H-p պ~��*S�=�_�y� �|�$r�[�|��0;�R0�d\�Րn&l0~��WFOǶ�N�����n6���-�mf�qN��H;�N$���|��=���?"���#{�Ӕ����K)}0IJ�>����M��Ȅy��V�E��Z^�m4�W�ww�����nU����6X�n�&���D���Ѵ}voto~�����([D�bA꠬��p��!��[+J�i��"_.{Y6u���.��\��a=HQ�Q5X��ցr���Z���}��j�V�ƈK��m�Qyqp[|7)���ⲛ��z��ߥ�w��d녌��MJd� ����D;)ӟ$`�!}ƈ4:������o�hH�1�H�Ēh�q�ȋ&�]�	���*z������̽9���R�ߔ(�H���s�gk�XS9�Q�Y�.1�Q�X�-��A�
S��
�i��o���o���"�I��`�"7��J��7��Њ�6n�~�I[���k<4,L�\��Vp��W!�Za�����j%)q�>�r�=�[�j��W/���%�Z��S�c?��z�.�ªAv���&� ��=���t������9�clcG!��mԥ�)���j@(W5[(�o)�(���3�Sb#���;��7�+Ѧ�׹����ZF�{Y��s�n�4�Ih>-P��'ԮІ3��Խ3�k�h�h�����.x" ����g�[E}-�#�*��bB�Ȍ�D4�kN�ؼ�['����F$�!�?Z��1wCr�e�[�]�XE�q��3��H(�m��&N��҄����X}����J,W�����׻�N�ϧl�ƒZ�����RfT�v���5�Kr݃e=`Bn�� �B%mu��rK#��y�J����Es�P��-훾ַY��g�4�8�g����be>8�}��d��m3��u�!���&��%��~�3]tot�ۦ*R1�KH�&$+>2ɰ���V��l c.ئP,�|��l��5��tK�#+�u�=a�:��	�{�S�WL� ��/1't���^d���v��Y���\g��i�e�<O�{C;-�(�*p�Y/bƷO�B�H���ل���E������ѥ�N{�tM��d�%ǣOa�WI�����"�����X*�΄O�����v��&Q):p�p��w���<o�����6FZ�M��[�V�m�B�qd*��hS��^n�M�@1D�y�e7����r���Jp�!�}�
�ӿ��.*�[=�{n(?+X@EdO�\��ԩǜZB�7��� Q��;��
V��;]R�5�FE��>yiQ��-���o��Y~�p��~�	{$ק��<���@ƌ��y⤃�ւ�������ge{v�5��u�ƽN��ޙʑ�`7�X-�};HS���Xݝ���w�@�zp*C[��jK ��L�P�^��0�<��y����j3S�����^2&�	�-�|cʘ�����Cu8hD�t�Oui�?����H��&7�h.�v���S�oj"�5�ZOx��O�[�wK$Z&gp=�Zҋ�`����x@�T~o��s&T�<jPM�Ynh�u�4�
�!>��;��9�R3-Mzh;"c���j�Wp�Nɀ�ra�C�qf�9�� �����mA��\�*at�̧��J�����|ka9��+"~���˽�)��COѮ�l�8[���(l��M�e�e��8��i�^i��z�p�� J�*�)���}�{��Q�¢פ��{M#p�,K��>���r���%��Iᣝ��s��T^1l�������Qhark��&��vBJ2�m���P$w'`��Й���5jF�{�'D^*�ڈ���K=_/%.�_�!���]Tv�2��ۭQg�> �Fnj)�({���R����,�b�l�;e�I�i�[ڦ;����{�B�cRiB$���{�Z
7����\�ޤ�Z��t�#l�$ؐ�Z
C	M��Hя�r�́b���p� �+ۅ�R)./���(c=�'�
��f������I�|���E\Hq���9EΏ���	��t
1���r�ΑF��|+׬y���Fo��t[�Ǡ�f��O����$�޵�g��K�1��1���E�Z�B��z��xtaU�	��!��eZ�����̝��_A�h���QL`W�Ke�0�s��K���5��?���w�$i}L =�������0�pA>V��V[!�fK��iD�d��UͷT�I�4y�a�G�`�s+�r��M}(M�)��9�n(A�,j~���,�pJ$�������8�l�p,��3����<������6�	�,P����r[�K�!R�7JjT�ͳ�?ːkn�:u���^YO�L,mҖ�UKM�Ȥ噗��߄������Lޖm;��
����%-�6�G��SF���u�5�H @��ofL�G���V����{�!��%|C\�o��z^ jNW��0������+Hg��zh.܉�e��HqF��������q�� ���~6]���P�Jc��+�v�c@�[�g��N/fI��{]��Z���s4ݢϖ�>i�:�X\dD�}��9�a�X3'\c��X=�����
�>3����䏄�C{�ֻM�@v���-��E<k���8D��U՝��%Lό�&�^yq��\JB}ÁM����sIcn:˴?�aW���}[7:�\8�y�u#�3J�9��^f��]}4z�t���/1u�N�f�ʺ��>=��{�0oz�kMY_�����)�f��Z���� �df�Y6�{Z&�J�a*?��8��e�&B��z�~�z�λ�<j�*}�s��c\뚡�$��f��ֳ���������l��{.%�x�e�p��ǽ���)��M	'r�*�Vqz�U��!æ������ i��m]��y�eELBs\�:0��)B�.�ԅ��.Yu�-���#ڪ��G����{/���Fؽ��w^���~7'N�#�YݍP�Uj��Z� ���c��kl�|g������5W'Z��|_7;'g�Mᢾ�a��S|�w�"_�2q��K��T��X�C&	TycPOv�*t��A��4`��K��_PQ�2�ߴ�-��liW{���|���b��6�D\��p}���ۇL�X��X�4w6��@�z��:9�?^�2P<&i7//W�%�[�ǉ��#W[����	!�s4"
�\����6�����e�����F }\�a����Å0:���'k�)Ӡ�E	�"��Bw���e0�ڽJ����?k�A��UYp\&��̬�gS��8f{^⹔tb��l�~4{?��;�k��O+��" ����/��)���/�	�\5p��o}�����۷� �X��{;B���&�_�Z��G�f��gLa�4;�<���r���L�t�I�^�n�M��q�=8@'�yc��aWF��ΫWG �{�X���
����Q�5!����I�c�A�=U07�u25Z���W��*)f�����@ Z��5��xۂ�g�`�6��-spz@j%#����%��%ð������
i�����yU A�j�:vd45x%���\��g^�����W�gC��n�--< �?�Н���h���5e���^���u���4�H��v����s�k��F�u�{��	z.O~ː�k*��MX�ܾ�1�����ؾ�T�EI�y)�23�T-�*	�:�e���O'Kތ��W d~��75	b��Q�H#�p��?���۸i�6A�`Iu*`{�|i�Vi����/;y�u��?B�.��c�m���I�8
D�'�����t�Us1G�7A��n.2�[-?v��6v�Q� ^���+�D��7�"#�۱�8e|5��'#��̦:�l�E�����2h�r=�a���t�o~?I������~X2�ᜑd"���H�������ͶjG��oFk*���g��tR�l�K>l�f���J���F�W݌�]]�>��GQ�W�t9]gI7�z@�9%Z�Z�ˁ@C������)!�f����B	X_5��ݤa���v���U3ܳ{n��+�1�?�.�%Gݐ��P:r�� u��|ju+%8�D�?P�=�J=������˷���4�B�|�>����	X��Z��+�&���`��y�e]�*گyO��[R��/�!	�Tj�������Kv{�vc�=>f�JW<�,x0���k�^\t��|&�`e������r���v2���e@�5� E�ĜzB��{O�#O<?ၹ$o��sݾ����ė׊�2�pD�FJ���`��z��%{ضb��ܠ��t���'ݣG}�&觮�H71��gg��@� 3�g��'�V>�@э������K���v�ƐP��.���N�ȩ���sc�
�6�U�v�����������l���@�8%������m�Jg�;x^� �-�3�.t�ݻ�1	X��h8k�]T��6��ܢ�U�����L]�ō`�o��%���R�z�cr(K������)
��
}(e(�[��u?z�����H��x%��s������/���NP��=�Q� ��ӧ�ܶ��((#�g*~�Q�\��B@ؽ��wI�V���e�
�9C��lE=!xj���gK�9T����xK����X��T3���WM<�<F��� 2%XP6@�;����M�F������\�o�=�
�i�r��6�F��/�WI�N���U8+��>�����������j�]EE�;��s�fcE�#��-�Ĥ�����%Q�V2�����;hL]%I�et͹������(Cת`��P���~���P'�:�P�v�|-b/��<d�q��Q���af��!N���:����g���a�UvzlRh�$�ւfSu��$�hof����D;��Yܬ�].v����ޭ�!L�]����h��[=߂������KeJ�
��0�>���AO���~���k+�$і.	�7���0h��;������OP�D��	�Q;�;��F����o������"���V���6{0~�<�.����]!�M�bԄY_�޴�w�!�����>�̚�D� 2���.�oy�NֵJ�?4�?�vr�~B���.z$r�n#��_�:�ROě��U_�f�H�XԉUTEҒawڦ��zm�۞a:���x��oY�p-�J/@��99~�ƥ�H�D����䊡�z�a)�E�{��64k֛)�Ǘ���#+\�c�XlJ-2����8�ȡ��WR�ܜa
�=�Q�⦏���1�,	�t�6Y�9,�)�tj�'���tV�e@�S�[��]6N�������Q�D]j\��
����v����ǥ
�����f�i%q
�=G9�0�M��:K�p�%��E��l�U��]�{���*�Ӏi�0Z��M��Jq��Q%)�,ީ&2'�����o��9�����1��6YXC��T�lO�X�n�j��x�_��GY��\���kK�(�K����ue9��G�s2����h��B���B���v<d)�υ�M\=q�4!�J +M�Tt8ڭ���e�S�Jî�XN�#���iY���D� �W�FA'8 ����bU�?�O��4�c�o���ƪ���|�J�\1 <�h��"!u�w�M�E��������4�{�/A6�7>���漍�i�x;���?��<�5`���B)i�,����ڜe�y�5�Y@ԡ3���b�d�PY��J�tlfdaK	�����ӗ�RX��hWo��P�.]��K�
�On���;qE�C�z��`�6ڊ�*|l���璄la�݊X���������8`\P:�����K���2�ma����g�07�#f�Ne���fmyn?u������
��7���! *��'�7k��U��y�V��>�~bB�r>�)��O��oA��9��1�KV)�[��"��,����#Q|�N�_�&j�ݑ̢���w��e�@=��ֳ"��cd/ ��<O��uU �9��/yٔĢ&�,;�g��ʘ�6��2����Coig�T�2�BX![;�a����׷�q�h���ê�b���o��K�e��?#s�Z�>Zd�)����|��d8��&c4<s����=T�AaIv׻��t8�L]X0,9���?&?] ��N������[`��y�v�M�g����S�My. *A���٣eb]_���S;�]P�ͬ�j����&�J'܆ ��οҿc�����P�r��e�p������M<��&�y��MB��/K3�!�ؠ��ALLXS�/3U�<� ��p]j����BC%u1��C���
�k �9H���;s
h�:��<z�x�&{�>t�w0|���>��g���	W�8aN��	Ef���f1*<]pzl��GI#���]d]�X���0�M��&�zO��m�������W0ws�N�������xS���H��G�H%x�v�?\vil��k*v�����R�澞*q��X�m���j�#�����}X� �:�$�M~�m���ik-&_�
�o�������Cζ�d�����`���ӽ��Cp�J\�HPCL�M�EҘz�a(�wh�ZT[�C�"�	<�����>��W�ŗ�N�OUi�(��١8��yIg����;F\��w�aY��R'����Oe�^��.Ylb����s{��_�~����*EƷ�1���V�@n��?��Y,2���#��y�?G�m ��49�-�q�ʍIZd�e56��3��撤�q] iUXj'һ�_ זj�(�95�>�Î�����]W%����W�5#�-k���#��=�`5��w#p������)�om��D����d��va����t �7珙-�x�^s���"��p����QtW��$�y�Sw�)��d�u���R��,����%u�<�Mn�f[A]g85�('m�q��K�=�$-8k����eQ �sn�%'�g0K�h3����C
�
��i��
�o�k纈�x�6z8~s���3�Y��HFB����v��o }7�k�*^�A�hZn~�-�)/GWH�9>�^�B(FU�KB:N�[� �r@��h,��\>Q:�i���"�4*u*թ��R�;S�H]ؕ�}��������aν�[
V畈SeMw
�wA{���r�F=�����>�9�L4K�q��(yuR���uM#��&+X��f��0��!��93�l^rK=����	�w��ų�.� ����� ;�K^v�]�/��+��xl����5�S�{�!ZO�$>?Ò�L�s��3t�S�[5K�~�rW���K'[I��BƯ�� r���̄�,)Ƅ!�L�Yq��^W6\�039K��ՒJ�D��袧��Ǒ���ǋ�q`U��r�����B�ݬ�N{��\|�Rp{n��������m�
�k�Ԕqd^����.㞊�x�(��F�ME�ـ����8��L��tV�[�w��7"�K�Jy���\��1ţ��{�J��YD�G�U�clw]���c(���	����ˬ���#�+��d�Vw��}:Y��,����j�(.	�H��$^=&��Uѥ|i ~`	����
v<_�#ܑfS�Y�����eV����G�(���+%�o�@��i�ss	���%p.���\�4��H���ѩO�{_
m@�J�dl����+ѯ%=�o�aY�,d��	�]�gi�D��ٮ������w.n��br�4!N�Z��x�g5~�6�c�4aΣs�-�@Hݭ���M���=�������i�����"ė���Y��5�F�grz��� ~�p���;�cU�o�� ����O5^^���K.L�:�`uxib2W
�O���h�	�Bj��}�����e @�D��!����X�]S�e��m��vG�\�/��:u4���gS�2~s[1�p���Ha�2������t��1�Ѵ�����s��SD�S�Mp�Om��<{k�Q����I�� [6�.�� ǟX���/�l/ �ᅖJ�3g�����u��ţ�����3�������>ڕ'�����<���cӝ5*�n�-�pQU��Y��'�a8�5��� >p[ ���3����w�6)��\j;���OF2z��ۏfCe���n�0*B�G�/����y��-%��ױr>��/=o9��6)�i�����KNx">�JtF��>�ml����a�T*�@z��츦���BR�"H���~U�O���=V��9����(�-�ӗw��_���B*B��j��!3��et�#�;c&r����@�f\~��,	���f7�f~�����] �y���B)�a� L�Yg$3�x-Ч�nV�\�۫2s�y���j���#���B�-�I���d��Η?��J'����F�K��y^�<��iB讵z���v��]�ah�*v�P�.e��p`,��YL���]��e��H�!��tι��M���J��\�b{K�7$<�?����+7��q���n���%��'�:+T_��-�Za���. ZBo¿���c��@�F��� -y�J�- ��
jE��>�Ǧm�	�M`j�T
V�'�����ܬ@rc O�fQBMiݠ�^-Y7��:"?�g<��☕X�Y)L��C�1���n��Cp6�O�_g���VP�?I�x5&ш�أEm����X��p$�{"��-�}+�L�N�\_�#��<�ܜ�h ����B���14f!��{J�VE�Yw@�D�Z��IX��(N��i���z�
Z�-U]{dϑ3����������������p�@��z�{=�����2��V�ψW\蟰�k���7>m��Iu!uN�^�H ��D7�χ���2������i��w��>s��t��U(ݐ�-�z�p�����z#��C���
eY��-1q��&�\ӵ�λZ��"��#�P��	.��fՍ��/��	�g�R.�z�����7�+&4������<������?g�JǷ_l[$����.H����|B�H �_�W$F�c@�����P�V��>������&��4o��K�Ƕ��=���z�0P;֤r~gJ����x��^���Ω�18�3�T���Cj��e�o��3�Y�J��+g�`֒
��j���3AA_k5��V�O_d�����+��QHc��:��KqxB�^�Pq�3 n+���r�����$�Xɾ�e&��J���[��}����Fd � �jy��YZ`���$%��;���h�Yu`"�ܱ� 
����A����E��]����}n��b�x"<�<����0�~�Cȼ��%0?=�N��Tq�Y���V�:�\�$��C(k ����adj,�n���|$�h���/Kv���I:���%6�lR � ]�	����|d�Ǜuӄbc�����*�(��(0)����8�ȼѷ+8�O?��J+y��e+��hA0,�:�ɯ��āq+*��U�ldw����a���<��~��Pܻ*{�`Ҫ�R�c�2��p�(5��W�G��wo�)��j�=g�TOqd;�}���bE��@�{����f��YM��7��&5�`V��T�U[bW�|���NP��QD�����ӱ!����lD����DE���{�����>��Ɇ�]�EK������n�=(�Je���[z�o܌!Vc���1̳Aˎ��W�\D&�Fj�ⓐ��"D@��{�<FjW��p��E3�A�2�?�A���dR��r��u���]t��-j|bl��C��!JR���`��^��3�0Z2qE��b���v�jg�Jv\�
y�q�o��kG��L&S�j�M�"夳�]��&��+0��3�ê���P@�Y-"X��$���oA���9g�=ь"��[I+7�uV.�bzfx���2�z�\�z*	�V糱)V�&��'1��.����0<C]5��oAAZ�MM`G�2pB��g�	/
�����r�^�+
�
�H�ԯ(R#ǏI`�~��`pu{��#6��<�H��W���()�"��Ue��ͮ:,F��Y��(. �8TN�f�G����p/�	���'�p���'#�'B�� ���b��N	�֭�Jt��'񐑥��������׬(B�n[�^pυHC;	��ˬ7֫z4�$�_��"�-��������?�ﲲzqu��M��t=u�JUo�nVg�O=R^QT��S�3�l[0<㲊-���W�Iv��H�>`
����"�
�Ո�)C䬎py�U�V����hO�b���O�.O��=�P^���!�������:x!G�;y�D ���e�� |�HK��g�挅�� h����&��D���d��d̦���	k?��cm֎2#����t{�I
��	a�6w`��Y.bbf�#�	%��|�-��������v��2r.9�=����^��QQ��w�ޯ����?.����9�i�_b9��v�u���/�G�]�z���ieR�!�"m"M[~��"F��#`�N���"Y^�t��BU���K�[h�X2�fGO�����Ea��"�*/z�B�[8��c�Qj%����G�1�/�l��,�HJ�����{�.⑘}�'�u�?�������&`W[�K���I���Q�*1���'5jM2���ٰ�����!��`��"��#4W0���TY�e�؍�y?d�FC�aߗ��"!r:�H	LU�Ci&
��&׈!|�ěCn^]w�"Y������5O�<�j���Ä&S�{�ݕ��(p�a��'�'NG�����Ok�{�U�w�]��
9����V�OB��Yx�n���Y�����a�i� `N��~��\-"���o�4]�á@�aJ�JoJ^�/�M��%�*,�cd�ߩ��!�25��9�Y�������$k�,9�$YG'��ҜX�*�L����o��G�R	�絅�FT��^]���g�*��k�ӣ��^�x���4ȅ ����v��5�c7ǡ��\��M)'_
:���1i���5�8ՠ�wﰴG����h��aGi'���VTnR�N��̢xBU;v8 �ꈪF���<qA|�F��
��C ���"\$V�DU1D�Ԭ5��#�Jz��7�q)��J��b�kl�EOЖ����:C�^1ۄ���H�"�n����$(��p?3Z�)���#���P�ez8T�n�c-XY�׿����#��k����(֢�f��������J5�ΰ���7q�Mm��6�6o�a/�[��S�q� 
��=��ͦC\ɓ��=�j�j��0-��k�8;�F��m��'qG�)��dw�T-�)x�����pW�.c�#��]ؑK�O�N$�-�.ۜ=�%#9�x�26��q6�N�x1�w:c���-)AP�U���j/�P�2�D��fMU  ђ�(aN?�dGu���4W�� γ|��o3�/.{5�7��|	��$���.nSN'QDiF��B&��|��9�/:67K�����!J�4t���u��7�V�=A��E����G�3VQPa��� Rv���~��3�L��x%k�b�r�/�ak�>e
X��9����u��/���k���9L�8'<�"���0�AEG
��i`���K,�K�;�i��ֻi+7��|�\R��Kz�1����+�y 8���S>�?����L	q*���>���.2�c;T�12���./FmO�󻻆�=�=�h6xH=�W��v����y+TM"&���/p2ݳ�@���fѤ�~�f����s$�zbv�  �+� ��-��6(��+����c$%%�4��CYB&��qG�Iu>.ӵ�f|��GԶ�������D)V�E�����Z�X
���\��kkZ`��3�eg�}�m�BN�b�6j���P�n���P�f�0��舣z�wٴ�9eL�z�k�D(�teJ��8_���k�z���M2��0���d��̦���xX����J�(�ˌM4����#G�,�M=��\ȵ �S-���r+���:�����}�I?��z�m�9��#;�ҽk��(E��А���"�Bf����;��&��Kb"6�/d����s�o���(�V�e��t���N��v���ϔF�
�)��;>�&�}s���?�S�u�/uaA�0�P�E<p�1��Y�g��yvr�N�`�UӁ�@��@H�6�ZƦ"*��̳v=�U��_��b�@'|ȳ�%y�Mz���v�0�ya�z�7u�k�����ы��T֠�?��n��>0h�O6ZtBp0�����oK�X�/��):T����y�7�M�$>��1A���+/�x��_X�K2%�+��l�/�ʩ�m�k����Z�q3�-�x�\������]T�G]����={I���U�ȬV����#`l�H�C��R;����V7���2�p҃7�č�+615�q��P,�$K_&�b7!���Gϙ���.�Ezn��^i�D<Ӱu�^ �\>�;<:t�P�D9 v��EdI�q�锇8��-�+��<����O����F"��6��Ӑ̧V
 Ps�t.�]a!��>�O\y�h=w�np���o�#����]\�r=�ZΜ�s2��M~k�����2�芖������_<��f��+6QGJ��¸�P��
�;��a��6B�A&2ʸ��֯���3g.@�H�y*`_p%�
{Ǻ�ΐ����7dr>�.)�:���I���Z�Ac?�ߠF0ρ�t��}5��(�
�����l_�M���۟��$I˛T�Jy�M	�W�r D�K�q&ξy	�\�	�;���z@��O����\�m.O��8���g�ױE�8����d�M#"�ݤ��KЏFX�y�U$8)rw�Q1�[�رI�=�Cm���VT\�W��IH	q����Z���RVOl9��tQ�+^�HB��1`��1��~6K���{kjpb�9In4	p~6>�O��d*e5d3�R.5g9��a�b�A]���u�@��*���3h�6$�0�n��yR3�[����_���.�4%	��@T�������ズX`���TUJ�\%/�P/�h�ſ��墰ww"�\�K*<N��"�C���jeӚ��"�I
�,�uB�=���]��m�v����(QP�d�Y28� ;��ҷ��A����dOG�-ꊵ�g��?�i�e"�2B"�&>w-�T�6O��EY% R��r�����U��qs�]�P�nw�|�0�޲ZT���ڙE��k�"F�_�~z��Gü6�b�	�jC6��G�Gu�\K��Kr�?.��6��dj=�W��3����h;�ZrJT��S0#��v.��$�0+�7<�*+	DaG,�w��Ծ��^;*)�o}��}�9�MD��{u:�������Z	��,��;͖���^Z���X�Z���C���Ү�R�����2+���lV%�oz�g߆!K!��v��sO�|�:D�QEVQ�D`s�j���Ƀ���;�cw�w�G�re�B֩T#�Q��\����õ��
�����΢j�h)��@�l ���8BQ�.욅*�aM�q�m�w�l��!�p�R�h�َ����l|6�Q�ȩ��-��Ml5s�����K�a"^W�e@lm�]���;+��W���`��{���z!�����t�Q�y��B8D ����h��ɢ�3SտAgh��~�h�x�O�aG,�/�,�>��!�k��ȼΞ�h�d�,ō�j@���a�_#$�龏�K)�!k'��u�; ϯ���.q��9��GY��Z��:\�|�"/q+�fh?���81h{=�qՓe�ÿ�N�H��ɓ�s���a=W0×�I����H�1c �:���T��ς� �Vr�
�!���1e������/��j�z�뷫��r⽇D�L8:�䂬��n� �v��>���3S��$D�&P�(w����9S�SU�c��Uv tdȧ"1u�����,D�U(nh���B�W�߬�F@��/D2ehI�<�#6��yƔ��K�Ƙ�Mj@j�s�'T�k3X{������'�'��+#������-�΍��F�Ro�DH�;:猞YbY��yN�,�u����vC��\DE`fsj������0����!��-� �e��?�w����ga�����<j�����u� 9�_{����_�UR�1�E�
[���:��Kd�uM�2�R$��W��,�o�c����\s�mY~�u�`M�K\��!˔�D��%1�&�w��sa��~~�R�Iˈ����E\%��R햘�2Կ�F.�ϊ@����H-$;�a���/T�f��Ui��Qu����z?u��J��z�����Y^0���.��)��̚ �K�]?�oG�ّ_n�&�O ��%�I����Ng	%b�(G�x���7��g�-{
��*�����UCQ���B�Ҙ/�r�?g��gvÍ�v����)eR�*S��,�?��,a�X����v�f�?z��گ��`�B��Ղ �Q
�0�I��ę"$/'P*(�����2ܷe���������)�S���`m.L�_�v[UX�%uT> ��>��6�ܶ>f��{��l!���'ǆWJb�;��(=�����-�l����X�oԌ�[`]�"B�;n\p�p�����y}����\���9���g7;��+�]�b�	��x<���1ibd�ԀD�ۆ.�q[-��)`�!�ɷ/�AEN�iKW�{d����$
 !�t�~8"ُ����ؤQ
� ���g���|�F�Qms����-�S�+;�(?s�����Ḯ/��ns0�L�o[d()���,��
PD�O@��������ʞ���G��~�3��	�Qb��l�}�+;���:�����߶���R���ڻ�G�{�b�B(H�#i4Q~�F�Ea�H\�`O�Rc��)�Xc�>gb󯍞+�� �h�f�q�Ҙ�EIH��I��w�4$A1D���#rؿ�&�� W5eʩz�xݰ!J9��>�[��.�[,d,��2{Qz�uF�仁àG�ιi*rk�A��.>�1��C)`q�;���yJ6
�����`�a+թ�S�G7���W��R�����jD7�pq{�k$u�^L��h�oz��6x�6A:�!�	�ȷ�R��ߢw���Iw^�P9����a�'Mp���"Wve��j`��(yv���+�=uT{R\��C-�?A�}X��g���u�6�"̛���U
�ۘ|�ضa���s蛻��, 3�g%{?��6A-��d�էi����B��bwe�_6f���R�߷��(�< �#�������è��zз������i��� �����^�[��0JJ$���±�b@O�A F'��y�D*��X-I9��j�Ja�W�P9G};=���P���n�!Ѷ�q�oz�w4���Dm i�������or���{�G��]^!���i��ɶ8��>��`L�@_ڲ��c�
���J/�,���+�g�Ǔ�3���V"N��6�=W(�ݘG���b�@70UIT�v�ްO����*��?�YwڟuYUP%��m,�6� ���B���Ka�Q��6k�dd�+>k�
��0?*�����#�CӦ��Z]#�Jn#�Z�����ow����7�� ��+�K�������?d�;��ꚳKҬLu;��,�^'�oU�S�e�}�P��^���l-�w�615KH���u����?g��Z.��Jo����
��	3���	���4&�7S��"�[4U��}4�ˬ�./�G��ͷ7�$�w���k��U�Uʏ׃���m�{1el�}�%Y?=.�ňˍ��nx��Z�Ñ����m;��c�:5��e�i��۸Ҧ�6+TP����ڴ_��x&���V���B�����q�J�1�䵦��H�M%�vO@R�8�_���ה�]`���Ω�){I�PoU�I62�pZ;Y޳���X��?bro�����d_��i���f���O1󅍭���г�U�!'f5x����,5Q)j�]�W�بd�ӽ	,��q�=ٰJ�B;�F��3��&��hM��B�7�ُ��KY��js��A��|vvΌ0�'���4���@^����[�xW���^7g�7���,G�Ӈ����r:O_M�.��'P#�Qb�5� �$p�K����N�3�
^)/i��4 �}g��S��J�/��"?I��R0fr�7d�_��ц��>,�0���JG)�h��=d�bY�r&R����H|m}���ڦG�� �W�ٶ'(ć
Q,ك��Y��nk�W����jJ��J�r�kI�_|=.�OhJR:����ǰif�ޜ�W�^�w
���X�A�Ì�4"=n�bEJ�M�ђO��Y�8o�]F�7�Af�����Y?Y�����,^���X���M�Σ&�	���h��~��t�[�%Fʍ�Pv6m�tL54_�6I���b�e��8 �����RMv8��(�Kp��:���I��9\�Ċ��?[z���<�:�_�g�f�!��$����yo3fVl~z~K��a��x2ņ�6��P�����	=��L׸V0߷xM������$W�������R�����l����55��,��$N|���d�#K�ƚb��s��$E�V9���!(J�"��A�s�1=�u �j�z��EZ^��g�T^��u�s�]=xC��BC�� 4��Dױ��^�����iR����-uc������ie����ѽ����'$��o��i��`j"�H���}�%ȿ~�j�Ě͠Z&'��~��k	�ŦՃ��鰐TKy�t�L'���%��zU�Ɋ��WZ���8l�iS��7*�����/X��>^��u�z�Ik���f&��s{ϣ��9�u<� ��)!�eD7j&�:g�<��W�~�V[�V����%��9� i�@�aWݰ�����O����������Wp�8�A;� v�G�.�Ub�.H�، ]�U]j�o���ߟ����i�Re^.�ح�z�}����2����u؄�UD_��*o�J�<X2�!���:��[PE<���%V�'�_ϣk��U򒧆W�DQ��~��zhG�'*�(�c%*�d��r��x���
F� }�c�`R��)k�!9"�mĢ><bi�|.%��bC/^$*��%��z0�?�Cpq.�]6�e��"N4B��8?U�&�i#���5��t�~VB{�3��q�:j�K�~����,@h�<��~�1+M}OP��������)S�v̵~���jw�?�C"��ڟ�����r�ՑV#��8FdY�C�Q���,�a��e��}��/gZ
7hq^ݱ�\KD��B��~�j��!��ܳC����D�}�w��� Uӟ�ufD[Oćк�m}�{E'4���	���s�F���ox-P�+��Ƽڪ���o��.Mʃ��$l	߲�`�E�1�ٮ�P�@eB\�RjaLwIrS�	[��Ho���Gi�������Z���Z��I���84�_�׶�i�,N
��%��}�`������
z�7����
�u s:~,�.� �~���܁{�i�Q���J�_�J*&hL,��i?
��fA�"N���0�W�|��d�����ˤR�p�E[� �F!˴��q��[��b0C$+�Icn���Q,�_Zs���Z�U���p��tC���z�9��8��R ˓�b�yW���������L�+�����?lUC���J빖����2�fM��w���LN2��H�a������)2�|�� -	#�Q�J����%YN&)�Ŭ�x�u��|��.�r��y���'�O�uSΛ�@&5��-�uW"�E]�o-����$W80�8��!uo��Vya���Q����w��CCe���{0��#���m��a&>ٖ}g�TC�ߟ��ߣ��WVka�$�Cv!���>��Vzr�qc��L�!�)@C��>�����fH�>��ؘW�6����r�눇_�X����k�gU!��i�7�EZv���o$�h����*l�c:YcD��'�]8h�>�#���:��'K�e��͵+��m1���!˄`���Z?�y.x-���JyZ78�y! ���5Ȟ|Y��. ���{@�[*��>�c�̵\����kH�k�	v��rN��[�;�3��do���o�#�ǹi/�&s��������{*��5��63M�k(��N���qVsX܉�I硺���Up: &^5���Na�X��p�<@�N���ֿ�0�/`1�֑�Ó���>��3��@�^T�8_�U3�\4�W�Dq��RG����h�� ��,_��f�=�ܷ۶�v:�!liB�8�N�y�+M5�!�hZ��(EM�ʃ�\0D���8  T���7��ҵ;�n��;��J���/�q�6Dc�OQZL�
Cc9u$L.�z�/{��\S	����m&����w0��s�Q׫c�Д��M��:��.�`����~y<���h�n�IQ�������1j5��ϴ3f7B9�'���(PtF<O/uYAP�22�A��S����tRi������LOM�������R%=S��09@H�Yp9�v%S�rrn?Z@�O)]�l�º�SaXf�,uZd���}�����ٛ�A��y�N��|Bβ�]�&�%���{�=V���Է�t����"Y#�o�}�bT��n��l��2�)�5��u�*���z��
cx#��~3�h��خ�,�w�5�%�"7�J�8
�/ܨ�d%�z��bg�ғF��HNzh/�4��5ڵߌ��*(������6 ���G$�am�L��H��02�t�Ho����-"��ބ��i�8]��%F���{�۹������A_}��@f���Z��0V95�a>�s���˹�� ��z6?��'�w�F.�>����, �ZC1��_���w����#p���[�H�P1��du<��g�70��$Ʈ���fx�v��7��������?51��jN�21�|����oma�� ��>%��Y(l�|�ʛ�9��/z��|L:��О)t��+{!qpڊ7�;q�>��YT��᧴([sb��������6;�/�is$_��2�t*�y�:�0[8���u}��S���n������׃rɈ'��j<��/�$m9�]��g�W��Vs�k�k��|	�� �##�&}�w5�O��kL�q��N�e�ػ���~��7Z��x�*�k���N��c�Vz��.E �ح����ue��1���u�������2m�|�׉���+�z�������M��l3�m�G�(Na��lKLa����H�c�My��M�0�*i��A����H��qg�\P�8���!%��R���
p#�Y ����&��+���������8���ō{���j�~�T3��,��bxyO<���.ns�gT�'����].�Ij01��[P/�6%8�]T�@��K]s���kx�d������}�o��!Drr���+h�2�̋�@�`e6�|-���&q�q6�#��t�8�:x����j3�.��?�e�������>�K��"H��G�ɒ�>�MZ1�[�s@�͒���+@��:����%~akDLi
�R�	��#)Uy�[t��~�p�$)��2�C�z�f$fW�Ր��x�M�a\��	�J��Ĩ�q������3��S�g�R9���r5�(��Љ9�F�r�I��&>���L[���.���[�FD7W��S�S[Y��g���J��r��͓:㖼�Dą��7���>a�(_������E��UJ�a��4��\�9������si>�~�����]g���	���/�SQ�GL=�B)&�"�����=*.�f[kH&�Ga^���0]�ZD,�ba�'��c���0���9m��.���~D�_[b9��l'�śB���Ľ��ӷ'W��E�PE[�mwy'VqgG���BI�	��?O��H3'ul�W��1�2Qx�L\*���o/#a���>tE��U���&���f��/���6W��;�Y�Hf�Y�_�tO3
�e	]81��op����;ґY�M���y�DMW�����(����M�n�[,�ǣ �pZ=q;�Y�О)�diE�q��7�_6�?��a =b3��e+�Ȳu&~�%2^��h"�ߺVd�m>a������o� ���<�Wa|���\����u։�q����|Gn�E�p2�Ñ��A�ի)�z�YgD����zyf��^-��&��<ք��������ۛՂBP��O	E��î��bvW"��y:��=#���b�	Q�&j�k��z0�ws뺈	��5��Lxf�E�F�i��{�:�xv�	c�n����U��ed�Rѓ�Ӝ爰��pfQ�BU���yl�g�=*����h���0?0�Q�0%J|�oUrG�B�T�uk{���&j,����O�	�z\���5C����%C|��
�k0+P�k��I�!��\+�I���>�U��H�`�$�"(e���0%��C3ًD	ޠ�M���,^�N��Y��4Z�7]=K����.�Z��Apr�h4q��W�%8w�yA����qJ#�C0���T*�[D�l������U�vh�Q��r��g��7Ne@?xv9y���h�{�dg�6Q�
����\����+xI�Eӛ��N[�2i0���!�}y����z*� 	����¬��4\��L�B�Dj*��<�}"z�CY��N~WU�c�������d'l��9�Y�4ه�3A�~u������e
�Sx)5�=�f�U���ӋWa�{v?Q�G˶<���x�|����t�N^�h˶��@�_�k�8�&���Q1����93Ȗq������$=�$�7&�O����\�r�H>�(&�bmص�"u}I�u�ѧ��c���b��罿��z�DL�o�w��Q���d�l�*��{��w�))P��9�&ٹ� ���n������\�G�h�AO3B����~Y2$�g� ��О12]��W���Ȯ|����b���#	"��8������F�����!�fM�i(��C�Fx��Ϙ"��
h�r�#��[[z���;���p �#�f��:�g\�G�87<���)P@�U4�J��B�h43]7l�����ov���$5��!#�s9��*��̛�hc�lT��V���*����_�E|��zrn�n`ϔ����Śg��ZĿQ�+k6,��_��)���5�V��s�r�8輥r��_�B�����+�C'�Ķ5G|uVr��o ?���X�o�b�����?x#��T�	P}�<Yʐ�]ֆ�-M�V>V��X���M�$Y��ɺѳf��4O^�@Ǡe��
����!S=�����t��+w<A&4��[�	�0�����Ic��Q��EvB�N�X��7#�?�042��+Ir��!Kv �bwNƣR^���ʗ�&k�&���#��$Н��=D����2��蒄�������pq�{��?��C\c����i҉��X	?o�܄\�/��Z
]Y�=p֫�O3㮪�{]^��	��P)�-<���F���ț��,v��a�����]��\`�"4~��`�	8�.򩯾B;�YC�l3���O����ָ�t*Z��|)r��Oa�d�i,���w��?�����E^1L�)����E(��Х�Y�n�]�DN��7�d��)�LE��V��c7@;;/�!��������@"(W��E��:��$@,��G&�`��.[�bl-Z�/U'���u��3�z�E��-�������$_C�	1��2�4����u^�o}Hc���e(jI<[��P������C�zE�GW���8�}"�U��l��H��A�GE���]v��ő�#�áN�CS���"*��@�	K����pp�X��U9�� �f���<��Om���Wږl[U�H����7Vs	��#�Yh�\��>�dq}f�m{�^yaZ����E�X�"l���r�D�0ދ ��.��룔y	������xW�-�7���5�[j-m���ɚ���Pٵ�L v�SG�U�2W��8�\l���J�*W��;�{Ԭ����øM��M{q��5,7���?!�p�E��͗�A�_3��o����=z���UG�B�AD۩2�;�~�e:HxA�P�_���CN`״�"M/��q��=C�t�G"Kj`1ܧ�XtFL��i��x�}m1J���s�
�,û]"�1!B��%� ���&5T��M��x��\qa�yWj��}uI{r���{{g_�k�'b����*�e���*=n�A:>0T�1�=I�L��8�O�:(�$1ȼ�U�-�����[�����w���dxR1l��A�8��v$l�|�{�@I��x�!v?xgr��ܖ�Mf�0�F��#�+0~�)\��R�Wyac4ǎ��:��C�ETFCB�1� ��J#��5QNݫR��m�׼5��>(ݹ���m����K�3�:�|n�Wt��˚��{*�s�Q��ƛ�Ԫ�.8�kG�ske�g�J�-���B`����y�}7OT?�# �K�f�,��'�V�����l;!���>�i�*~];�����vs�>%P80-&m��ɜ$�F���+�A��I��W�b�2�&X�b��������[yAioi�c��yx�L���y 5�#<��vF�"�ǖ����d�3XG�9f���F����"�2�Lz�ye8[5�`�� ��SmΈ^���+��(A�%ŻjB�y���j���!^Zv�|<K�����E0���}I5���	~ɦ���z��(q��'J.�Fm�la�b���}#�:��GVj��r��H�@��
󙣕�;>�:vU8M�(`ɔ�䐟/�������*�gjJJ�E>�Q �H$��F��}��|���qgKm79��k�d�3ʰP������w86�^��G���k"v��EV�7������͟�1�a.݀H��8���`��X��ns;bGT3(�%✁��X�C�6{v�����+�yu�]/�X���Nwo�ث�ˤ�����/�d(0-���+"h���Xu��f�ގv&��2���|k��F�����7��h Xݬ���4�Q�ni�7������%E�oF��S��&q�ċE���Y��o��}�p���z^�
2cU����c[$p7��N���
rϗ���O�)I�a�u>�fnUe���$W �!#���y}��#زL-X����睒\�W�wPb:��V�{q�0p�~�EI�?��(�9�!Zp"�H��D_�P[i�3��r%1�=?ɽj��U-F
�M����ꓑ,��mk�bT�(� P�N �8�l���ZbȜ3������)X��ϝ��6SV�)����}�B�����Yx�5�U��HR��(@A���}�Z7Y����;�ذox���m�Qx�B	$�3֭���$Dv�;\��fYX��Lf�����v���򱸴{z�b���h�"���[)���^<�\.�s�(��˝A���f9{G��X��эl|�Y��4��0	65���S�W��h��f����k}���^�D�iQp�����/��_@���I�F����Ym�3�����k�D������j��b�=�?�����EQGۅ~e�Ѓl�(�s�˱�F�>nW�*#3������R�#�`@�����H?n܀���8v����Ǟъ�[/�?������@��%&Ŗl�d��N��=��;���,jC�GGuM�����f�2̼�LQ��,GQK(��f^ϋ�)�ѹp[���Zg�);�s%�ǐҙ�ƕ{����ו5Ԅ�
��J�����N�ϝ�i�W��^�ux����%S�W�sC�a�x��tNH1L�n�B���uOz� �_��f�y,��6]i�:�Vx���i��P<�	Ѩ��Q;H�0��f����k�LC�*�?x��J񅐞��H��R����T�]�&���^/�;���qV��1R�}߱D���C2r,O\�f)ދj�4?�|�ۣ�쏅҃�G�����K/d~X�l�������֡ K7po#e��Щ�'���b�@8}`���9Ѣ��|s�c�E~ ֊Ez4*u�(��Z�;|�aּ�N{��No�*� +�(xb�#:6�M�>;"���_+j��Y�N<l^�f�5 �aOPX&�)Q-J���1�scUB�)»�sc@Y,���0A!c7���z���<j���m�|b.��T䥁���||�{g���h��<YH���}�އQ��S�����u�@���U� ~��.?�z�ΝA����]r��/�����*M���YK�I�Z�b�UE���j�
��m�қ@���|�*f�D��h��2˯�4d8A���V��@�\O�2���^F]���_"��ަ`��u��YA;�|�-�Ӓc�YY��Ig���JN���;E1OZ�}kSc@?��Ԣ�e	 Y񪡋;vX�x:���/Ɨm���.�fo�!19�e�#/��hf��70>��GIoCx���W��j]���F�aY����O�٣�H��^�삏�7W�'��F�.^΢����b�붫X)ƴ^
� �L�Z�t�3/�WV^�dz��p~���XWp�ҦS�7T�~̜@Ocj��Փ���㓘uhe�����Zh7���V�������x��1�q����w��tQt`���Z!f�9���Ӧ�����g�\[��gI�1h�Ƒ@�e�K��)6'�yjs�p>S!�������F�?*����d؂�P|��2SY��"jN&!�n��(B� � ����epo8h>d��Z�&�zg����D�k����U�!��2\]m�"�nw�~�]}�s_�GƻcX_���Mq�I��Wa������d��=޸��#��fU�����aM=���9�oT�N�AFAo����D��Mi,JV>��A��L�fҰ�\��G�#o�}�X��"������+�o��6��r�
��X�%he|�_O�N1���T}��g�3�D�G��B�?���w��E��ͥ�I��%����)u!P�;��`n�:t��%B�����u�>ه�X�ا�@�?�K�ɚ~Hs�T_S�3��,�bX.C����*S���-v=���V���Z����
�Ub0� Ks�����w��m��6����^�0Q�Cϔi�"m�#���jߦ�3u�]�o<Fa��(��A�޳���R�9���)�WIp�f5�	�zβfjJ�|FM��� �N�3yh�.Z�P�d����9�Wy�w {!#��UC,w���JR�f��'"1��1m�X��`������<��6	� @����w���z�b�-!o����Z���o���耰���`��p�B�SW����h(w,b�(B�L�6��Kw��Ǚ'��8���o<'��Hx[/�6^����27�� ��R�D�0��	�o33�r���
	闤[��@�;��6>�h�2*����ś��"ۮi�
��u���_ݙ������u�;��Zo��l�.�"�O$��K�<>�/k��l�tڼ>Q����h1udLdgrtEV?���9�9�8~�a�zr�G [��x�%�,@fl��P�ٴ%M�[$��NK�`�m t��ic�ݰ
��z]ѷ�9�3ZB"L�Yh����I��"ͨ�#Y��=��DI�����7M�U�{*�	�yO�GA�^���c�܉��b'O�޺n �PVx�ɏW��W`������U+cz��	�0y�~cz��T�R�[��/T�4���I�-1�6�~����mirF!@�j��a���+�����G�r*+�0�dU
�9ÿY�(�����3o}�_΅�zZ�I�3&,-	������������e2��Z/&��Tzmj�Z���<�R�-αu��XxQ��~\	D>�%��t{�x�z8ubb&L��s��w1���U��w#;`v��	x����H���2H�BK9� j)��Z��B&�[E-�N<��m���Psl$���D��6���Pg��Ȇ���2�����6��ݓ�l����[R��+���`4��F�>�۷T��\Q�rh11]�d^4a��0�(�ā�E� �*��Č��r�s.$��&��T�z�a�ϡ�A� �5�B�?�|������C=�Ԉ �p`4ݱ�M�o��5!nĭ�9�,qd�N;!F�o�D3��.|TI4��yh;Yk�Q	!XN=6Q�t��n��uDϼ�_&�ص��lU�ι2�����5��I'��A,��J��/��r�.��:�v���b=���p"�����x� k���Ы�'qb{�Ur8�O!ʿ$c��H�"�D���&tK��o������%hvd�D&���n��"dͭ���m"�k�Cߑ0�p�ߝ�:��lt��z5-[i�f8�n������DK8.�Rh�(ڙJ�`: 7�v�.������'�K����{f���uX'5��W�du�����Q|i��4��Ʋ����J�0:�p�	-a�����ozg��ئ�'F�5i�������*.�S� �m�<�Y�>YF|�I�2���ﺷ(���i�L���Zق>��C�s����HJ��dYhv�_)o8k���Q�Z��9�x�ש�r�����	<�q�<���S&,�Qin���SE�O����rq���xm��4HF�A<���P���E*e l5~����G>�C���Z��6�[�����_Pw)G�����/�3��s�辥�Ҍ`�2{P�y1ֵ��酸�G�����'N��󁛏3 �Ù$^��J�"e�
5}P�F��eK�����u���X�����i#�Z��<|/�4���yfŢO�)�$û-?^l ����N��0�w��&{�pV������Y�^Y��v��;�v�M��?Y�3W�k�?�|_lU\��Ŝ��r�5��֫����jP�Z��B��YnL�S��hc�TN�GJ�@� �3"�6�{����U�m(llB�FW�[���vmxT/��Ο�3Oa�ש?�9��R�<�u����>h�-��"�u�r�/�nbox(0A�n��_K缨���zwe��+�)�1�kZN�����FZ)��wZ�z���6m��ˇrA1�L�I��a3qZ��'K*��z�[W>?��m�sSՄ�60wG�h!X�c*o��b���K�R~8�G6���ӬmDb�ύ���'�Ӡ��%cqQ�Mޱ�c���C�z����3�7K��+����f0�B7�a�D-�e:)f�b���5���@��xA�k������\�FAY�s 3}n.���I�.���I<��,��D���y�·,-`h��V���m�����ĳó�E�4�e5�/��:�5�5p�c�M�������@�\5��1�|pq�6��$��e�Pq�*V��c>��}<��L+h��0�'��1�Xհ>��ς�A�PrW��!.�g���C�la�\�"��
h��Y�z��d�q��́N�O�1�"���`}q�;�jY0.g���ڙֿ�r!9sĄo3�lLf�ߊj~�w\_�G(���>�0��,S�O�2�t�vI�L���C�gf)U��;aw\����{?�X=|�zפ��5�u#�ݲu���RZGI�o|�� ���0e�w�T�`Q�q�s�P:���JD�'E5��W�H<9�٤�r�Y��^u%x;���;O��P�r�(�|��p�����!�=�9#��SK�i��?�\pE/u)�^�2��"^���iтu?������^䂘A� !@����6�l�n냡��6�6`'f{��T4ݵp��KDϦɖv.M�@�-X�%t�܇l�as�����X��Qw�k?�ߛҳ��j���J����(s��Zk���-�"�5�[s4���t'/��(�qku��	�p­��H��|�9��(�r��^��A�Q���4���Rs}�@{���P���������C݄�H�J�_O�?�] k�lATڐ�����%3m� le�w����C'�%ai%5�q'u_�Ǽa�wto>1�'��.��{�xV�f�Og��t~I�K�]b����\᥹-��Ӭo�4=^��|�̴T��5��R�8�7Xg�d��~	��0Y�~z�Ρ��Ϧ����@^n���o�ͯ�J$���N��y����#�K���4m�0�>��WP�f�9����ZM�,#_��4ƊP<4ا>"����9�R�]��b�\���a��B�b�]�ˑGa�G��)��Ӽ4%O�	̧GCD*�{Ag�ӎ^��	ز�<�G0�D3Ch3������cȀM�#}��`�9`́�7�|Jn��UW�+��<7-y3Q��Nu�c�H x�u8�5}u�o���o���BK�!�Wm[n��~'{�7S�qw���mZ���Q�q̳cA�jQ�,c�5�HO�b�\��6��0H���#3]��`r_u�+�A_�d��k�8�dZ_��YJ�oR� ���8���K{���3�7���Z��z�g�� �8w�:�8<k
�Y�:����*7���1%Q���D9���^�=zH��s��*������I��ޚGw� ha5_2~4PH��:~unc�ɘ�ag��S�Mr��zoc�)���C<����Ņ��D�6-���l䲇G�B"�)!�@�'BB���r��� ��g�jr�y����#I䊤v.�.��[g���?�ۋ�������B���0�� B�x�?�%Nڱ��FLߧ _<�V���}��1)s8M<KC���"�\V�?"s�=� z	L���,[ٵ}_�ԡ�Fn�n�fh�2�זL�s+�S�ة��Wڍ׈0=�T�%��'���H���w�8nJ��W$%Q��i�ɇ��2  p�r�����ad_{W��z?���U��D)�SqeW��r�(Eb^AR-2���E��x*�Bk+#(�� �&�9��d����om�]y�<�6���Q�K��+{��L�Y�Z>-�Y�(chk�!G��[]3��1��h��䡌)pZz�G�>9L��๟��#pB�*n�Z+�?��O� 6���D�t�B�� "��o����`$�F�;Q�����A�/��u;��{)��i�@�c�U��ҡSЕ�����7�SG࿤�uA��{����,�&�1D��4��ۘ����x0�癯���2��0�Y_2Ew�Έ7� ��IĜ����E�b0a��4{�0���]��8{�oo�Ҟ+��&�{BC����-j,�I���A��g�|u�bh�-P�[�/oV�'�+s�}U79��/k������;�wyv/�dYEU��@[��uz�Є"<����Q�7�k�tN��|G"�|tp�,~�5�ݵ�,?
-��N9�C�D�B�@��-�O�7)�L2�洠����=�.��G�/�?|˲-���Ze�R'7�޷Y�Ih�H�hݱ���^��`p"�мqa7Ȉ	��p�J�5��(C�)C�~}N<��z��_G����W��*Mq���������!��Q�?�u�T��6�����z9\9i8� AX�d�n��6km����#����R�֟� �%c~��B]�O�a@f�~�+��_f�b�a��ǧ
�M�e7���x�W�y�Q�8��XT-=7饆U����<G	�zT,"���F9^�������>�:�K/�#�ũ�cqn���A1��m�'�q�1 O%{O���]��CHbi��{��-s�P�~����n�$M�$��M��g�������W��9 ��WOu��aG�	��7#��ZS��}������P��g�N���+W������v�yN`��%ϻ��E`yܻ�,� (*#$^���a\y����v�X.ջ����+j9:(�e{�%�̰��^�F�̓oJ���i����j��n�K�%٨�T�4��vFWM�����yGyb�@�3k�0
	[0���Q�����a�iß�wQs��8� ޳��b$�{W�Q�[m�T'����hߋHM�kcC�ۅ=(����.7^�o$\ķ��6x�@�ֵЂ��B������i�F�r8�@�*����f0�8LA8� ���*K���=�R IgDQ5�$(ٓI�s�_��Ѝ&��b��׺KID ?C�&蘼
�C<<SJ��ZN�f;��j�Z0Ė@�v}f8<�z��! ������(zo�U�M�8 ����ed�U}3삌.�*�-�8��'O�!)Q��{ۡ$��������׋�l����CHT�,1i���&�A�u�C��� �=����c"�����li�:���k}�Z��	���)���ܑ�9j�%ZnQ��"��1������b��J��I.m}�u������U�����[��"�^z���ki!���lw��1�r��٣Z�ȐO��N?������=�,'���#�Nt���L������,��8G�ɾx��Bb���g�o$��ڇ�q�'\����Ċ��|��AJp����D�fw�F��!:� j�"������A����Rg���`�i�|�8M��sk?*:�����I�	�TG����4#�� ���M/Bo�q�ȴR���������+�y�
���}EP���A���^��^��8�mCg�����b��ξz��;V�7��1�~��^�HL��^w*n�	.����c�>w^�H.����7!�x�%�i?U>�y�(1t8��O.��wVL�}�M�����&��_ZLV�p�X�":,x-��;�8��p��#"1��g$�ύ��h��9���tE�HP�9�l��MϘ��y7��CajxQ�r&�H\a�%�7z�C��\��;��x�(�I7��d� ���4I��f?�Լ\�*:���W�|9h1g�%pݤ��Sfs4�DB/~}ݷ}8J۞�s�����������)
<�u�U��xQWs�)�Ol�6�O׵����>��XA��l��w�:� �t��� ����d��N�ad΢��w1A��z�MԈMé5b���׼��xeNKl
R�|��w�o�j�\_��K�����Y�����x�|X�A���S�	{j�~o�b�`��NT1{��]LK�FC/6ma�5�����AX���j��o��/<u�1�ޅG˂��{�����I��p]�����������;a��s���7x�#NCB�p��m`{��+��q�5�(��\/a�؆�[wj��d�t�����F�(�8jv�%��Q�ڜ��qN6���s.���ߞe2�;I��Q, �� ��<�a�&����Nq��|�=,�ǲ���$!�l�#��
�8�uim�5Yl�p(��4�ґo��₇�'	�稷a�ӑ�_U'�����%�4X��3�}2#o�Eȯ��0ΙJd�W�S��X��5�:]�2�xY
��a!������u�D�t�x3����T��Ku�X�!l<��)��,|��k|���_�҄��Z�xf��ee��g"�ԑI�t="�׺�tG��ă��&��و1v+)��Ll�@�"i2�~�G��߆]�K%��������ݍ��8q,�b���Yِd+��4�S>�����J^�l\j(`�����Dz|i�j*�w��+M�媔��K�������`�.�~\+��"Y��$
+[`8�g U~s8�����0�����t҄Z��42!M)�����2A���HS�<�_���N��}�U�#k�wO��?Fٚ��b��m�]J(="�=���;,�y�1�xg��ԑ]ٞ��C�	K{��U@�B*�we�m��V ������F	���گC�pY��ʡ�or:�͔ �!1���*�@�s�j���
AFgFm�|�	�n�LU�Ot��95K��~��o�;���ū���Nw6'�u�0N=��\���;��GXmit�fl�QJ��ō����ҍ����F���رM7�[�:��bu@�7�=���|";DR8&�凿ka���H��[:��H�Hk*�<D����-�����i�d|� �EO�dQ��l�m2㹮�l���k���d�����z���`�v��$7+3��t�(�+��!z�G!���(��"Z�����8�[�_Gɻ������ɘP>� |���:��w4�c��[�21=���j����<ĬK�vm��.��u)�J�����gAҳ��'c�s#��|-�7��>(�������]9� ��<�Fª�u�Λ9a�+��K��qJ��H�q�1�C���u���{�6�{}�|H���t��L#ʛ��1�	��c6{B`HI�j�8l�&���Vic
��8H��1?[T��i�`�r�|��ھ��+
�����Rz��K��������. 6�%��B;�	<pZ޼C:k 'Wa�P �Ÿ��킱���3��s���Fɫ���j�zl�%aۅ�g��?�>s��_'N]N7r>x)�擃�V:h}ؔ\���=M��̱sI�q ��vK�Dof*�>��n���D���}��ku��p�9Z�XJg�a���@�b�t��Qq�^O��w�^J���p<��N`G�o�<�ֱ����t;�m�y�!���s�E��j}C����`��/�r]`T����<�HZ���]
l}�
�إ��T�"���&�<ܚ�Ȧ����=���IHk`��s����,)��`���)���_FZ���b�-b��B�w_��-w�σe�#X�ƒъ��T��9�ʘF�"�^���{���N+����xKp�l����,�{"��r)�]��#Il��T�e6���N�ʾ���ɡel��Roԯ;��eME� �Z">�DS�7)�uX�����^��sva��ce@�LS���9��VO�?\��g�߭7
Z؛clc!���ЊU��P}Ĉ�;����+`(@�x�O��t~��@I�t�6�;fM�a���j*ey<�ԐZ��
cd��[�;�4���-_�I�n\ΉNqr|1:���ؖ��<p);��K.˱�9�F{�� �t����.�_��s�.�b&�q�~G}�5��;V�����2T�|8��p������$K.�.J�w��J1ۄat�9v��>p�-��~0?�r�"�J_���c|���l�RD���U�%)���0�b-5Ĺ���㍼�m�R�8��Ѻ
0<���HXV<>�}�Ԝ�'�8���+)��?�8mMГ��\�#RW�4�#8��o)[�T7��(|ޠ���%}A������V�|Ӱ<%�I@H�F�t*X*�]�)���i�O��qcq j����OX�a����P~W̔Z��);���։��F`���=��?��t�v�z\�"G��:��(��	��at%�Ö��-MW1�{$~AÃr�p�Ih���y%"�$I�)V#�t���Ղ� c���^]��#si�<�]�; ��YQ|��@6��*���VGe���e6�\�F�C�a�\G�nSz�,�J�d�i���n����l�#�Q�䍠L��$��_�*E��G�lQ��`5��z2�K���c��1w�!1v�r�'E��"Е�_��ɦ�eBtD�����B˩��	��,@�嚆KQ�l�� �Y�s�i�àFV�Ь �C��cgI��}����K�?,��P=�`
ؘ�]q]b6�˸��u�J��ga ��m�cU��8a�s>]>��$r�N�p.��Sμ�����y\�vS/��З���-t��.�P�ε���q�Ӓ�l�_`K�ɭ� �u��{,IvC�Gp6�� �����v�W��������ڿX@B�{]�og�uu���..�Kmq�8s�{]e��"#vR����p�Ҿ�G�_2�|�c�P�H���;6��'�('�h1�w�����1%�����Z@C���b�����_���7�W<�"c��9{����J�o%����.R�"�,#}�k�U\����z���`Ԡ��ܒ�	p�!���:�
{;U٣D29H��^�,������n�z}�����S�"�u�{���	n��B��Šb�A����
�\��bB��=�Ӣ�r��Ú��>�G�I���.Y���p�A�cV�H_V��(���%�H�&]���,�Vb8�v 70�_���_�Y��v��)nF슶pK6q�62��@%O���\�!#u���_��l^�y5��O����� �tr,�������@��7{��3�W>E�?r'�[�J�S���	�b�!0�8�]��!��t����78�M:K*�T=�/�b�SLj�yg%tJC�X��<L��K����A�g�g��@�!v��/{�As?'ήs .Q����q�]���6e���4�G&�hw���x;�[#�����:�������'p�E���hj�bОYL�L�U��D���gW<�F�M��d�M��j +��kѲ��l;�/۹"&���2�tp~5�,!^<T�b �3�ыw�D�ӌ�H�ߞ��'�v[��6�� �q���(�/ʤ��7~̢�j��1��;Г0#�5j%^�<��;R�r]��ނf�n�p�A��?���#u BIO�����a�f-����ׯ��T������	n:�L�m�H�'�Y.��̧�X���Pv,E���T���T����L�D��뽳��;,Q��ȳpMH� �釅m�Ga/��x��=���]O)�������?B}M�����s��d��O�����o�Re$�IPf�"����c1� v]�,�8�Q���C@7���_~���3Xӣ�*4 �ٔb��ʷ�^  U��^.J� �
:��`�ry���!7���#@,�/m�3�B���7�c҂d^_���@�Sh7��q����cd�: >"·��Ͱ�Z��+�����⦬�W<P��R��3�T>����"^@�tݧ���X�Q���al{\�ͿZϪ����H��L���I�s��%�V�MsBR�#[}Y�h�{�KN�Uw�eK{+���,;0��l �/si��R�5շ���{w���`��m�V������'��~�,d�c:��ئƗ�	�p{��p�d�`�g�slAh�����1?��a�Λ�m�Yl?�"tHhd6BTJS�r�p��>�-�M�Pr� k��?�� 7�~�7 �脟"N���^�H^�Fq������s$��#ž�gLn����Qu��.h���|l@`�z���,�Sj�5��5�a8)��������la�SU��kR��;�Z�7ꟊl��v����1l�`64�68�n��d��~։U��H�7��A�4�zV�n^hT1QF,Eo�8"��[d����,��g��|��������q�̜j"ϛ�bF!V�RMe�Z�Rv�4�(���\})�{���gD9����SOü���ӿފ��>�*����>r��-	���5�U[p�P���pg!��py���Y&K��#�bܙ��V�lW�4rLwv���m�_�q[*�ź:��+0���o�r�����·3%l�1((����eo&�X�U���ub�A�A�Ho�����
���J��f��B\&�%��O�(V�{�]7���:�*���F������*1tN�2�J��˧�끹f�V?w/���;����|$�U1�����k]����`[�*�u�n�[�c@�~/����&��HY�	L r�����e�S�v]ݨ ;�������]�le/uk�ɻ}̍��s��
k�Um �\��X��b�Iߺ��1�>1��$,'�/��P��I�_o���t��:�M����}��v�7bh����Q�ɚ��t��V&r?�X%�1"6F,�͈7�7�$vN@���d�nȂ�	�)�Oy:Pd�#���4D��r��A)c�fMp	9ue�a�P\���4���U"�j��("p����ri�	� U?<�X�VF@xpHdB�_��zL�$H�Qm (���~zr��H��w~��}_ن���܅���`�X�r��*Lliz{
!�siB���݌[����a��@��Ⱦ����xI�)~�n$C2o���>��i����j��1-O{�ͧ�pP�x��*ʓ�z1�~W���y��0���/�hZ0'�(V��YT=�]y�)�O�;KۍSM4S�/ŮEu�v/��/�CN��Ɗ��~�Պky���6u�kVP��e��]�5S��#��}�Pm�v$�����=��W�Q����\�P헵��e��|h��Z�y��^��7�,u�`��f��N�W�2�lM:_&Ab�P�j��wA7ך�gpyT�؟��n]3s
�oo`ڮ��	�9��d�ɦ��^���e=��[i�[�rvH̗�'m�~uC������5�	�L&>Ei٠d�h�	�kl6��#�~K<��!DG��a�DᏔ��R�G@�{��j��,>9��l�jׇV��v�\���ZT�ϨC�g�4�&7(�|�	�yv���2�I�RVϦ��f�6@q��X7�_jm�}s�`�
��S�."��\����\l�CR���j�k�)	ʽՉj�@����}�ke�Fq��T��H$���Y�7��/��Vg�1������E�<1df��e �뼡��JL ���7r9�_M[~#r*������`�+y-����,J-f�j�'&T�����$��\����_�Oݦ�?,I�� �����V�:�m���,�����+/&Q�,���:�K�^�D�����0���d�O4��ۚ�T���X�ylp�BҲ�Mj�����HҨ�`|�`��V�{��!�S�|��;�L+B��N���2v)f"	�c�g{��m0�x'��'�rn��Ө|�
Es0�5���Og�B"�cA�MP�j���ٖ_.�@�����DIʏ�O�C"��nĪ-�G�i���Ǆ�5����f����.��Y�(��_�{���U���`u�[����@�[U�tpN�B�2���ZVp����M� ��������
u��Wo�V��B�T�硋0��sd�ze�ջ�w���#n��)��TŰ+ՁX}"~ �*�_��$��P��*E��ʤ4�������I�hHs�A6S�\�v5�?]®�M4���("����}G��H����ޗ�N��=��3���@���,��>v�D�=���kmp���Vq�-_�^~�V���=r9�@Q�}�H�����/>�딧P(�.�}^Hߐ�5�e��zX:3�e�Ef" -b�ˬ���U3P<	S�oOV{�k`~_%�P ;M���������J��vY�� m��C�eJ0��_LxMq��%�:�A_"��5�G�x�WU#/�TMp:�C�(Ga6�\%�Z���{��6��T�z�${��ǝ4�j�����j(����nQ�/�"��19�?$Sk"#�d~���P	}5F���U'�<)��I�#}��Ŭ��uX�{��g�K�z�bA�)0�%�C�)���wLP��QJb[���v��'|0-@�q��+kS�=q�k����{�R��Ҍ��|5�����-�N�l+<QH�%	��A�3�e�oc�Y�,�3��6V9����w���S��P̓
Yi���N��ȯ^ ���^�P>��e�m���i�ɄvW��6�_7�z�-��� 7@��7_]_��~8AD-��Y+�����VV_�X�i��;�`f�(qG"�i�7���kq$��)�tйe������u!J�~�d�6Ŭl$>sݴ8���|Ůi����}	�P���4���	��)2#B6·�ΊRfK�We#�活�v��K�.$ ��9	��S�xW,��m���\�O8�~�Z�����؎�C�QT�ѡ�[�'~�<Oԏ{���(G�7���_iŭU���/H�%�v���$ϔ�`3:Պ\�}�mh���/��di�A�F�~�F�`������ ��ueɊ��LS���/��y^�p�~e�� *k>\��5j�� B�䀝e�z�>����h��7�����]1�/H�g ��8���_��,�4�����BDW�x��6��TWQ�M"V���ڲQ�0�~�Pc�ɫ�WDY ��?�՟�/�3ݪ�]���+j?NgͿ0����&ч4~v����D��r�:�Z)�nG�C�fT��ʅ5�.�iADK!�%a/w�O�2�Gw�'%s��4�/�0�
���z��Y#e��Ұ c]��ͫ{�+�
�"�� ��q���|JM~ۦ��۞��'8y~�z
\.�3���bT�8Jj�z��O���u�?�(�ƛ�T^@Й�ٽ^������G��I߾`���"Gc���h����סN��J�B��˴�����@�-g5eu����dz����� �Fc�ˍ��;����>��Z�%�>�F*sO�}��u���IN��%{���1�k�ǧ�1'YN 2�4.�k��*]���_�hwGٙѽ�{���Մ����%��ūb����eAh��e��b~���td;I?�=�څҧ>0���: �>�%)�&dJi��~��R���L��]t�Ƙ�ڶ������R��Îlv4��]�n�����?'�� f�7�#����{δe]�
F���3��>���h(�/Ͱ���=}x�AJ�gM���2��3���Ga���/�֕D[%�-�.�o��l_hʛi��y5�\��#x�>�����K,-�&�/e/��¹�m������{�������l_ l�E��H�1ԟ�C�H%����&����9�O��'�}��ÐУ��%q�Gq�:�;3�5j�����QO"4ޏ�o[R#	�r���k�n��硴��@H��}
(�lR�~Nē<.ȏNy����~B#Ht��9�n�Ov�"w�5�7p���wha��2;뎠�;k��W��
��D��d��7=\�]�S0r�f�o�DK*�ؗm ����UD�!-������i7���s�u�)���@"������Ċ�h!xS�����z�W#X,��c����W��uG	���8���
�p҂����8���Ll�u���[*�\Z`Qѕ2ʛͽ	��N�L��o�M˵��#��_7����!DY�{�w����"X�����DqV��� 7��vi\0�۽gz�踱֨�X]�B����vg�� zlE\4{j/�.S�������c���{��<'NuOpఎ]�\w�T[���`��܄�xO���������/�4Ȣ�ܛ5ۺ��\�!�-���W�V
�@6�X�jOܹbarް����%�ᾕ�j�6Ϭ�"S�Fp���{: 5iWQ�F��.�d[��;6Hp��<MMF�Xa����"p��o�H s�x�N��t����`.P��)�����4��G�С{+(���=*o�(n�\�KQ�!,�vQ����OwD��e�G(�Y���P��ݤ�иj��J��y�T��:���q���� l�6���g-3��NO>��~�i���[���oZ�sY��@�M������4 <��d0�k_��EW�Mj������l��-=:yq����V\J^�\��XnK�ϒ8v̳�#�mb�t��Y�`�Cby9r{��G ��ʀ�A���mDt�j���c9��V���C�	��᪡NN?�4g�����f~(l����L��.�r�m�dT��$���L���2�� TA�+�Lo2���D<yQ_�H�c��.YY��&⵹���oG�t]�l��|�K$�d�j>[^�Lu*	��o!��Tw^����4d��?�.U~����7Ϩ��)��5�Ѥg�NJ��c� #����sD��l��Q�{�$I�/���K��7�=q��V�d�Ħzؕi��Z'.R�>y�ND9�7$K�a��$+|�JI3��ۋ�&Ż�г�T:1P�q^�l���Ϙ�4j@hv�^ -k{��5��2yۇ�q8���D��/Jh�� � {�B4̏��~_��i��9��9Jn9"��Te�3����=��#\������0�-}Q �h@����u����Āa�@"��耪l�w��kP�$|��77�Ӥ�[��$t��ꨌz�_�N���P�)�a��wmf��ϣ��Jt"�&�'��e����q��.n=�����/BS���^�V]o��w��zY4ZB�#�QS��.����$�S�3-�T��}�)k�{i>HG>z�u�O��49O�,Sp���	f0
�z+�? U>JvF���Ѓ9�н'9�P��Ĩ�S}^~X,!d��)�f�&U�~/�h@��jG�F%�,�R��Y�_A��B#�n�c5PV����ξZ~c��P.ϣaL�� ���A�M�t����D��A'(��n��tVn����PÔ^�eD��� b^,�����E���S�C�(˼ ��R�4��Z�����FŨm` ��-hާ/VN"NHx���Pm����(oƽ�� �Zl�)����!X.�zo�X�>`� ��zr碰C���Uxc���կ�9Q��WX6��;�P��Tl��"����]ݑ�+W�\�B�v+���潝F����p��?<��K�K�r����iP�P���DD�K�N#F4�R*���rN�l�X�����8��;ڥ�jo�2�f(��� �߂�3$���Ф&���1�6{�^xj�k�����M��ז��J$Ң����>�_�즨�S�%��f���}Xf��kݛYi�ʢ������/�_!��!H���4~�&j����-�1�6 �=�˺�a�ċw�~'[���;R4�,�3ǌ{J����6��q��ND�[�g�ܟ�9(����ugN��dW1�1q���D���O�-��*��X(��fT_���|L�?ܽ�p�-=�+ySg�_�m_��m��){t��w��:��pO4Ԃ��f�Y��_={��0(l�5A{��'u�gqE�y���{�1Q��>������O��o�Y�z�.!"R�Sl\�ҌzZ������ �W����+�|$={t/�Y��+:��[�1�NYC��Λ���v@��n��.�	���<uRX�l���K��`5���fૢ�:�-�X�2O���n
Rݬ�m�@[�>�&�5AC���Q~</v;���6����r�=�7�PX��{�XSr���TnU�Bq=x���Zh��8��hX@������טl(������_L6�t�h^w��������B� 5��8�u�R���1��0r7h�sz:l�ݺa������F��R/��'� ��s|�9yl��Ƅ.��uA������J���ކ��ȓ��@X�	�J�H��Fۥ�@Mv�'/��PgC8�ڠ�x/l���ZS���5��z��WF������2�wG|F��|�F����H4��,��v%E��O:��g���gO|���A��S�@Sw�Ђ��jB�<V8�]Y�$n�-C���M�6�!f�.��Z_����RyF�4��,̪Inj������>1��}!�y��`Zf�〈E��D��\̻$��=��X�cs�
�[>}٫B�(%uّklV��e�͢�ӛ2�pk䊡@�"~��u��L[Z귛C��RM��FEL��6�� �KF��5l�c�1��1o7�E�ajXu�!i�d�{�Z��!&l�6��V�8\����Qk��<+*q�����^�lIC-�VSH�� ��4O� !;��=��\�W�2��lQ�5m���x����~ܖ���lȴLm�݂� �S>i�������i����	s��o�����$����kO����_�ޗUp�s��Pѭ��1� DNB��,�4Ss>2�Tl=�J��~�p`PNPM�^��`�q��ڢ����d�K<�����|C�����ht�1�Em����bf�>as�):�2� ��U�7���`��d�O"��H40ݹ'�u\�H��k�U�o��t���J��1H;ˎӉ y^���b�+��e.������怋�퉊��-�����Ϟ�����j��2�y ���9T�v�gbi�^|TN��U9w"��]�.�p���l,&�|gB�󘁃5�*���|تDF1�NH�뀖�g'z�kzW�fBL����t��W��$_��}��%���L�B1���i�:�E��<�d�������왽/��ܘWA��Q<F�E6ß�.s����F�$�Q�^��
?�y����T��a�X�������¿��6�"�Rv~%'N��Ш�E����K	"�����E�������J�_p�JG�ʘ��!��>��Ń��E`�}���{���H�S䕟D��`!�Ͷ?w�������3�����O��G�^:�f'�X&>2�E{SH�����P�)6�@G�A���:iu9��d�k�E�՘8�?��[L3����6N�>=]x���.h�yjazƱ����>>b!�s8Q�|[$�Q].C�>�J����������En������x�_q
0�B�C��!���9=-��%w�<ˎ�Q<~�>�f�(����9ĊK��y^Z�L)��=G��?z�T�ɯ�������F�-���|M2��Bʇ�"v����H�/ϳ�Y��"���H�F�	����cqs������~��(�iOyR^�/<I��(3���+[�4+8)�	~39�-C<�%sB��j� ~R����W�A�e�|,�`��Y_O�=a�S�et�a��I� w��{o�B	�x29��gμ��'N2&C�Vq�L�� �xч�E3��󥺖w�"���E�l���4�zS��H�"
��z�*Ai�e{^k],��P�
Y�|�L���<";�9�2׳ÃK&V5  Õ��V����;���l����6v\y�p�x;
��VS�O$��lx��L��� 1�/\��8�_��̤���o���'�D�u|D;�q�C"џ�V��F���rqt�W����Jw���H�El4�N���?Q�尕Їsj�c!]w���~(T�^�V��w��'B��ǭ����С�d��
],H��@J̍�!#Y+�h��V@F���nIy�;�3K����a��$�	B]�G!w���;n�L6~���`�o|/u��Ә��{Ѽ�]^�[�((�&�I�tw,]�������y뢯r6_]��.� 79����ѻ�w�X�&�8�2�QI�~֠v\Z�:�L�L�1M.��J6b~*$XJ��~��7�P����NB��kE��#�3�����!��q�y}�8e�q1~���Ӯ����"���`��� G&y[&�9������K�8m��{%��]fmr*UN1�S���4�}����m�V�oG �/���8�A��]7���k��T^�����)��sO�����~|��d�]q�w=�ǻ�s�As'q`���mDB��/�ҹ�eӧ��yx q3�l^�>��#�����6�wR� �\���4|��3B��voJ9{_�����[y�{��M��II����|
M���>��9>���Q�*��Ek���O��X��+I��h��^��P���3v�-��Oe�B����=D�k	��G�$'��)��~�`�a^��ǫ�S��L\c�v�D��nߙ�Ǝ���G� �z����� �
�Uk�N	���)#$���RM�2��`kLtj7�ήm������ޟ}�q�cR����6�F<�8��tћ�9"�_�c��I�½�e3쿰M�u��#�����dݐ9Ԝ��%�!qq���̳���(�i���]���3������1�
���WV?S�#�[�K�^�|c��-hZ�{�3"�MEr&� �)��|����4j0�s]nQ���8I[yӕ~�,�'6��t�`���kr���G�N+�<&�hX֛�J��g��;��x�[5ay%�BpTg_!��M�3�H�X8�O���;{ӥ��I"�R<��)��P��:LȪ9�9:��f��*q�:�#�/آ��*���2��^�淵x��X�'������{��I�m�4����3���bV����g��)� VR�]�vӈ�	�V7���<y��Լ����t�K�g�+pnҗP��Iå6]8�}�����2s1������-��:M�I��,g��.`��P� �xM��p�5�v]��_��3��D<�{���MFIp��ߺ�����e�C��w�����ZH:6c��g�q��&l�	���svľ~��8����*,�Zx��M����Yvy4���	������
f�0j�~D�L��� ������zٚ�љNFӘB��k�ʘW�y���J�1�g6O�������|W�5�,��h�d
{��v��� ̭�������U
�qo�82�^�ŵW2���mk�]�M����k���T\�4�{��e�aAq��&��n�����~$���e�BI?�|K�s���j��l8ȑ��D=�G�
�Uˆt�3���P�V��X�ؿ䢋=@�:�-������7	�@���QL�y���ʐ�'�|9∰@$��S��BuQJ���;Tķos@�,��u+�Yۭ)0bRsL,(�5>H�QF�*��U�v/=G�h��LP͒F<�x���g?��E�Å���w:a��Q2L������	���d|83�W~S�����O}}�q�Sr����e�?�G'�̘�=�P�r�����(o�f�����B]4�>��`(׌�.���_'uc���� ��G���	�ޞ�|C��������YA�Ƥ;>�] Bޏ!xm,!�cE,9~ �U"=,{�\�k���VI mdpS���u�� �;�0L�J���/(S�Xv�e�5�E�� �z�2�T�!X�h��&�B{_��aV����������e���	��xUR)+o9<C���n!���7�Ѐ[:nސ�����i���e����˸���E�d���o1q����)��>���
�i��r^�(\�����=�Vs]M9�z<���<�ϑGD�$��^��Q�Cy_��{�r0
*��OU���:!�x�m����S��d{	d��:û@����L��3+2�X����%���A�)l��FK�����&�D�ܜ���+����
o��H[��4t �6�Z�Bd�m�&�Pr͙���D��G.C�
��3�ȴ@��9�Ʃ,�����"ŕ8dl�- ��s�i#&��`���i[�NXoe�61�ؼ9�L,��o�t45�]8`h�$s#�a$�a�BǷ��J�Dj�(���4��R�)D0���m1��QL���1*}Q'��dv���0[
S���R�p�R$���~��q�Δy�T�.���?T�K��\#�(���Ѫ��2,��@�:����fy낔ml�$X��4i�g!>9��䐎ع� ڟ|��?>��<2M��8�J��*T%�O�>g�EE��p��Te� ���������|DCC8w�k��š,�5t�\@���dy��Σ���~M�~C*��U�Hq��{�+O&7NŖ`�p���Ҵ��)��%r��C��I�����*���S�qe	�g���i0 ��ɧQ��u�|���~®VLp��6z���^ɘ�}����еo��Ɓ@7��O�N��n�.�[��d~+�SB�$����Gq���-��$�����2{�xV@1��X�"W=���/yP��U��D��_r��`��7m�jOل<	�����mʮ���/����y�8�]:w�bV�� %cc��y,A��y-~��F�[�ݗYc��[����5��c����z�ϙ����i�ql�̀�����ɥY{�������ݬ�;v�D��93�*[����V�h5��q_���s� ���x~=(^�?�=x�� ����O�'��=J� E<�f�V����Q��5¶%�:?Oq�u*ʙc�il灷���l?O�G�[�m��֜�s�UsZ'�[����R���)���|[$?4����� ���,	�y�|/!v���[�*�nU�S��}u���ޏ�#cKy�}C�]���1���Ì���� �L�T��\v(XDq�v
�,�7]�������ގ�<g�$�I�%t�x6N��g�:n��>�y�MS���O��6�W�Ӆ���NB@�63B�$: ���)%�-*q�����0�9a� ڣ/��G�����g�z���4��P�����5�XB�n���
�F)��&Y>���muP�b�AZx5���	���K�����<�	?LT��2ѥ��8�Z���?G/�׃5� ��kW��g��*�)�gt�E��pg)Z���C��*p�R�&��5��#��Ww]�˛�7n�	��[��V��]���aM�j1o��<�:�M"?eu�B�FiM��$Jh�~
�%�X}D�f(�!�>�f��&}/�y%��Ǖ�ڇ�E܉
nT�K�8���*>N�6:�d(ݴr ���6Q}
l*�$Y\
~��9� j��S��)�E2~ �.2����'h
��g ���<����Z�ny�����PI8�R�
�O5��?3�N���M����	K�
Ē��,��FO��яl�_c��B,��j� �YE�k}2���@F'�( ���� n�k���g%d��r���X�K��M�#X�Ǐ�|cB��\V.�9��<������a�8KO��0���K�`:���� �/ݩG��/�S��7ū�cj��ӠЊ����1�Z���Kc�\@�����o��m���l�0�͑�Q��/�:uZ�X�PO����M����F�ϣr�ǎ� = YD��O�?+�sG&e�Aw���kt�,�`}^qH�~���)$2��`b&K���K�}�
/SL�T�0������a�1��s3W�����9 �쁓*| /2�;g��_�+R@E�p��1��0�����LT��sød��n��6��&Z�9�����@`�|v[�4�Mq&�Տ{��O/!Be�X�+�`��G�5"�d�A���<�_�B�>�t��e��wI�yc����z�L(��5���U޷Сu ��G����/��o�|��z���,�
l��9w��5B�e��:<4�n+�����Xu�Ց��N���?~-�y=��H>�!"y����@Y(OQS3z��e��)@�����QHZV���bd*��Ţ��鈹���)��A���%���1���`�N�w��7EҠ T���|�z|y���͸R&����������%�;���O�L���a�A#�1��}�w������6Xo�y_�@o�������?�?�XU����&'��b|=�3�ל.'y�Yf�\�$���
�5f@9hV�v��~A,��v��)���� H�	��=��Bb�N���~����^jD�^�H@��ύ�q�kt�ş�}��T����p�m��rv�3�Nrwl;O���g�ި��R�[o��O$�RR"��n�8��+^�9�n��j>Ț\�]�}p8R�'��c�o��
����r @.QfhQI֝M,�t�?3�=V�������ܚ�'.���Z��#~ C>��f�_��`�m2��!q�w�+�y��)�K�!� z�ē�+bäJ��!��3�:��ZH���Z�}��G��w���t0�3|{��B�Ep��9����?�9h����l���)ȿ�B���w���:k.˺ϓk=�'��N:q��Bd�m�W�D�� �n�Ց������h����:ɚ�[$�������?p�e��r������<h��F��9h%��iz���Ր�4YqL<,.1�?���Sx�Q1���)�*1�O��s�3H0*��-Z�8`>
f���3g���#���g��n9~>�ڎ򠌊[.w���Yw�I�����O�����j�V/��ݝ�FtCy~n����eeGT�(A��Ü5�]Č.\?7"Jd3�n��?�Ne�v�恤۰��-�)?��k��\f��cL�����爹J���x���?�:���gom|����!PC���d��Q�V"yoz�C��bE��V����k8dI�I�.���nRUħ����:ݨڈ����l]!���g�q�}3j��K�p)ˉ~��HQ眰�x�����l��|3���!N�O9�?�?C�d��uI-�E�]"���*�O� '=62?.j$3'a��O�������j��w��J<qo�̹BH�?x�8�������*<�y�.�d��B�.��9HW���A��.���lGpN��"��Zx���@��f��=���,�0enfm�Dú0��l��n�M��zjd��)��(����@��ʵ  U��f��!�@wr	_�\�_a	7���O^�(����+�N��(�,��XF� �q�NH��K�K���C2����_-�GD�ojN0��Ծ |M�WR)Cbj �{�˷#S��/�tD�Ġ���I���&m�F�R�ы 94^�r�*�[夌��+�DZ�)���uɾ�:� ���y�y9�D%�Z�NY^�qb�B��Ɋ;�J�xexwɭ�.������`㹀R��T+?Q���3�m��2���(|_��Xb_V�. �nt�E6��-C�/_�0�ak���Q����]0�'�����Ho�
�ڣ�)m����Gi����]�d����g.u�4Eb�t�[f;��PI�C�iH3�@�3��d/]�X�'��0��O�Dk�v��� �M�.7��[ȋեD���i� X�;d�����*\,>B�^:1Ŗ�%ei��R����ũ~�V5^�Ӏ�C�P�g�{ì���Dr>>��:��-�1�L�{ܔڀ���t�?�ta&@��8H��	���T¯�M�F�>�o��T�м ��I|��b�W�O��	�scmX�]?D��u.��;�l�xª&
b��=�[x3��W�@n}@���BT�1O�V~�?Ic�h���66������.���(��s%,&ȶ_��q�.�]b��4��Α�M�Ѝ�n�}�|���{N{pN�|[�N��Q���/Q��y�́��9%�:� ���d�'�o��P]�\��(�N/���r�tY�Ooݠ���*����/ᦚ@,aU�T���z3FI!���ϰ���@F_�Z>3[٢Z��MH��k���9�*.;��e������@h��%mhj�{��| �;����:J�����t%\h��퀜$��ʌ-�2sh���@XWS%����U0C���02�b�{nT�8��'������D�F�YB�i��gX�[�H9��|l�d��/��3g��`�Пq�!�&�ȁ�"2AXkZf��ij����F�jl.��\��^���LUc�云���?d���;EB�ت�L���`��@�A�nA���P磋�qx3�c��"�X�B;�X:������:�4�Z1_ W�����ϕh�)�T1Y�N^���]���*9 eP����]�f�ܺ�S=��^�	^��=�7��������������2���[��n����f�+?�C���c�E��z6�g��k� ���g�/�J+�Vb���X�^S��=�������]��Cu�3U���f��o�)�enE������	9㔩��(j*o�f�Em�u��-:yo�7us+���0-�a��M*M�Y|U\�a,��3��m��y��#���'o��O�1\��Dfp��ܸ���+�Ι��o8Of���%�9�ĵ��@�y�8��9*�eB �K��R�[�:��
�p:i�[sU�?���?�|3#ɗy��ݩ�H�O�������׀�t��<�X�5j���>kz	�Zz� P�FJ���%�ns`G���8�t��^蔜0��
��饦��������h��wx�����5nb	�Y1,Y��$�Y�S������%���4�u������H�Á��Z;��qT���?���a����ۨf���K��}�Y@�������?��ѡ��(���qPI�����4T�/����xD)/,� ���{*o���A ��3���9�����2+C��� �;���.�@�ݕھN�m����+�2����n_�*ڃ�#�̲�뵦�C����J=�!���'�,����H�k�A�iC�ǦX�]�x��^��1z7�ev�ښ��m&~k�Kd> p�Æ����u�H�|(�����}�pOʮN� �f�4�Y0p�Z�
IWf�Ƅ�=�zT?�|+\��2s�J�2�M�HO)��� ����V6>�c$�)���q}��S��&cI:�V�Q	����1 s��~��C�ǁ˛�'������?�Um�M����ITf�)����m�t���
�]�h��y������\8
:�[�n�'���v�հJ��.T�'���_���S��
���t�
p��p0�(Ԩgě%�&�ӌ��Zy����d��X����!�ciY��'�A�E�ָ-ox�z�L1v�Jj�"��ǓH�E����>���[.o%���x.y.Bx�EJUx�,�V��mj�-�Q<,��[ۼ��<$5sЀ��%�pQ~ZQKx��](nMx�F�ɥ���`���úU��X?�������0�2�@W���	�߭����c�r��%�TW,ȩ/�T���ŵ�f\�g=nG0�cK<[z��wc�}�99��}�#�P!�����Ԗk�@8�5����X�������8����f5�I����å��_PI��Xٯ �
�����re�ҭ�@��?p�`�.��U�NI�{��X������]��gIMIX�d\�x��(%�1���-7�CBC�WW6g�����}�W	��58�Y1�
%�/0�,�/��a�ɴ�!5 �{Ly�޵u%6Y���Pۛ�s빳�r�3���5��34)V�uK��u��g��������B�%+�s�6r&��;��PW�#O+�n�*t���^R�S�W���`�k>\�x�~B.��5!)�A��>���!��p�6������h��Tܛ[�o?ZrD�x[!HR��.�0�-��]�b�(6�����ef�2m�Ց�$��AQB�v^&��yX��j%�%5ܢ�vQ��_Cʤ�볉��v\IJ�
03��Q8�ь$��3��^��<� �������0�Y��gCȻ"�����xb�P{b�'�!X?�Uϐ��e�EW]fm"��ʁGPlĝ�5�نeMW
��4�JU�t)��k���39�8��8��T(1��A����Gu:|���xO2��6,!������{9�|P�{��OUM�x5�to��2�ޫ�úr��3��1v���{Pi���!���uy����>�MD��v�ơR�qx�C�?������RyS��n���P��L!���#"߇3 0�!N��ɻ�p����Ei����Ɓ�Q}�O)pC�T*CS��,�dPKF��e�z����H�֍_b���nK��@wu��v�*=����O"�=|�� c�] �ؖ�~����wݟBr����$齈�^��ŏ�~ۅ��l`q4�vHa�Q2��tK&�T6l���-��dd~D��/z?��wl��ND}��'���8w�<��3MPf�K�@��0AxV��� ��_���'��^��W@��D�<d�>Z���QOt�s�Y6&��P��;�=r<=�;ru��;�|��ӫP�5�[z4>���9g'��`81~@H`ܣH�4?i�,$�����7x�A/���r5U^����H޹�l�z攅�a���s���U���CY�{�� e� I3�k��G=��&���N����HY�\�w�'ђ�`P�V:i���Mi*�2�I낄c �U�HJ���Xւ��2-��X��V4ʖ��PCU�o�$A5�<Z����h��Vׇ=h�e�ީ�H	L�S%KY�j\Y������Kh�_0ϵ�? l�s,���yP���V���4�b��R�������rI���N:�w�h���~l�"�q�R�Y@�v��	��7Z6�rN��p�O=�tW��X�&�9���O�}�}'1@2�竨�$%�]�����d���	� ,RxO�=e\�F/:Q�j@5n�����K����eС�a���Z�Hhf�K�W]h�7;�n��/��T��쐖���F��$��5��6�mڕ����:�iK:vɧ[����������"��S)7~雴���J�5��r�Uk�6��X�趋Z´�y1!B�,��Z�үϝ��\e�������7����5�>h��v��-㙂4�i����d�ajVZM�"�\�}]lPi��B�G%DP �d�?@*z���A�n�6UL��mף"X������H��m)<(���NÇ��&M
��)�u����|.�j��:����{�����[�9>�O��M�|�޺�hȢ1`��w#��&&�s�ۜ`�[���s�g�Y	�k�^B����<O10��5N�2C��EXR�s��%e��R�Y����Ή�����A�{���� �k���q��螸��=ē��ҏ�0�\�Ñ��,�k�a1O�jTz���KsŘ�%����ԇ�r=C�y�%\��#K�<R�9���%J��/aУ��\Ft��Sh�>���I-ic��M75�W&���G��@Z?Y���u�������"��u�C�x<����pX�A�p�u�����_��QK56��˸��%#_Kp�CJSo-��*����ܱ��X�vu����Cu9݁�$¬�u�a�d�j��U�-|��[��P ���'P>9 S�9�Ӯ7Z��\�Q"�N�>�����_�~�;�V�3�Bf�%R]�K�����jO>��o�p�9[�]�����J��5mV��ƨ,߿Y���a���g��*�<\{9�AU���7NKX���s�fl��uZ+�\��௧�_���X1k⸽�	��A��O������h�	,���C�PY	s+��Tx��z�*�J �g8��z���v^���0���ɺm�8�3'�#�ϫ!��$����=W��$8�<�2��d��Aʓ(Z��5�CN�sQ�r�?i�O����;����!�y���e+Ёvs,�g�#pgR�/�r��9��Ё�j�N�R�_�%�=��f��˙�2�4��mn��p3��S�?FOr�������$��ԹO����~x�J2�c���+tM�fP	����N���4𦮚P���*#l��R&Mer�9��(�h�bǡC^G>�{�\�%�Hˤ�.q�ىx��-�r�]3�['	��C@�46�b.��pz@��ہ��GWg-�\��u�%���S���N���0 �x푁�5ÏL��^ �����+����~��	ޖ�� ,
�7�n��K5(�������1LVjￋ� ���.,���M�P���˙�m��V��W�&;����=��v��1�.�?ȝ~�tJ��8���y^t�>:�Ьk�H����L�퇪"\���[X�b	�-�8*4tu����Lzq��	åh񂨚��5ކ����֏���,���M� �z�$�ts�>揵9j��	��n�S�&_h�)������^���b�!(�V�����,����h�K�i�2uNR龬�Ƞ�	�J���=ٗ)��'�c�'�A}�(I�����,XUڹ��qePU��~L�n�}���%��64�o��+�6E���k�7ig+�c�ifi�Y�g��NG��h����p��x��i��JF8�r��CowP��<�5�Y�$z2�2����P���'S>�-V	���#�<G��"�q<]�J�l�ǺS7�*�������8��G�06$��)�����0z�Q�oc��8�~����Hϫ.&!0�~��D�����* ����r����M��6�K�s����xm��ތWR�=�j)mH�k��*I浘$���o�8��ׁ�{=x�|�w3�Wmx�!x5�XG��*Fbx���<�n���a\��겘4<�>u�9�9�Ndu��̹���t� |�J!o�y_PO��F�R��ʲI��ru�!*����h ��C�hΊ����d���8^6��w�O�[��U����E����gKjn�]��-�\u�zJ��2�C�!s�kS�U�)�	0�tW7�8(�-�M�i��6Z�w�Z��~����� ��\�A"��@aP�HgM��:�y��o1��,iy�����p�"��n:t�����Z�>���`��5)�yp�88����19��{k�?�����'�魯���LR����J��#bK�MNa_ s��&]�6�WA!�K��n@�ʯ������ײ��#0������Ӎ�着��ćI��m���3i�t�m~ʀU.��*�P�o�rn�;�Y[�`*��S���h^�
����񟎛n8�����n��]M�/LN�"��I�?�߽C˯��ϝ�� ~���q6��d1�J�0�2���㳎���ER[�pY5���H��$�td��~��}*�ǔ�s�>�x�����\��I�����)���²s���䡐@"�m�FWM vi�v$���3��4�ā��V�/��aT�����[�ة��]�ZP�p��ԃ�<���,���t�J@�JX!�L��Io��d�RV�4�㵫�a�Wt����l�^f����������)���O�Qx΋rhw\�dP��`�j��冩ۗne�ڰ
R]� E�=gK��z�� } �>����Գ��A���A��[�NjN���H���$��&_�`����g?��s �����m-�Y�y�'+��>5�����J��F&�q��{?�AL��]8J��M|�������W�o�G2�5�4P3O��?:��,��Fi~�(�벳�[F����Sz��x�ZF��G�"��KZ娋U'((�^3�U�o�|�4�������#�r3Ϗú�z���q�}�]�z��� ����ޭ�CZ9K�ӗ*�s0�b�ߢ{g���`5?�G���T�1U�T��$�� $��ە�2k���EO��9�d��1���j���y�_\�&;ڻzL��H�qmO��^B��G��DAOsg�=�E��W*Ģ�\O��>�L�
!M��Nv-�5X��^�M�ԯ�Ҁ�V(�#���x���(���e��nR���f���T�f^�2��1�Jmn[�
�-B�~�ț�(lEP��^�e@W�%l=0s�]��+L�;��_��pղ}�r�v�km�N���F)�찆�����K!��xو\�%W�3.��Pָ��?�[q���m��H�~I\��n��>ŋ�Y�����b�0X�jLyw���\{Az��7���C�0��]pn��3/#�s��|�g�h�P�Q��=oXu]�]6 oh�]R�eƑ���d��뚏�j�dH�}�J�$HjPopǵ��!�������߯�ƞq����� ���k��ڳjT�������ܨ���Evz��Ni�]�3�6��d6U�����-߷O�/u��<I�T�ڴ�� ?s�����W�1Ϋ����K<#��U�S�fi�E�~0_��	�D5H)�����;T�SN���V�	e�Tp<ާ$��8POl����[��	�Hw�t7�پ��@"?���:��ȈFU�Q*���Y�c��'�_��}]�8|��~s]d���}�n|S"ihV*�<q�[k���&83atF�S�\(Z�d���ʕX��G���Q� ־��������^QihX�=���p<�k���c�m�������R�$N��+��Q6Ǌ������,,Y1a]Qm�G���uآ��4|�9�N�����f%�$��/��� L��@�'�h-S0u8=.=nY������s+ُ�\Z��i<�t�,<�9��[= �
l�֮�Ԁ��y���G��n�����ڟ��HH�Y���;��<�Q�u�,�I�L��BH�W�g�j��E�����1Ц��,�?jQ��xJ��7s~,8��:�|�F^���d�bQt�ɕ_5�LM���P���qa�1�I66H4P���7�*V��}��Vr�+}�� �,��nD6dȴ�J־�W���u{�/�.�-��
�=ئ}���K�f{�U�x�~
c�7��U��2ch������qN�&��鿎$�EVj��H9U��N��
4mBU%|(��#۵ *RHG���-��Q��𢦓sO0����W3�������¯҈�g�9ĩZ�?�'��dߢkD�.$�@ab��ͥ>�)oZ��70�� �тV�6�"���"�ї����f�D&��8L1���h&Q����������ނ���J��@.U�$RŃJ�ʘ*���uכ�"�B��Z ocD�d2�v�7��M����$C*�`��5���}T�H]Q�s~������ܫ���f�h؇CFY2��=���%$'�J,��ʴG�ٱ)<�ԁh��\���޽��*�^�嬪�����^�x�|�w����N���($�ӛD���-Bȍ+c��V���c��3$����w���(pFE��-�˄��B���,Έ�)��b�hKz28K�-� },�&�D|"uc�)�E�
����KV�<�<�m,�q�{�컼|�,4f�� 1��y;�~h�u� ��(|rh��,P��\�˪"j�^�ض�&^�����I���ưaq�=�b�@�Mɦ:̉5��G��iu�Syp������B,|J6拎ٿ���z���pc�ad�H����10��iթ7�k�f�z���;]\�����-ú�"ElV��~��ϵe��Q��'�Ĩj�,g��P��J!Q��z/������4���S��:q@� ş�<�qy��L�x{Ň�īZDJO#�Y>w�|*I:�9s�Ƶ�^ͩ���
6�#⦄�sk,�2�8�`��{m�=�p2�N����<7!��&ڃ��q�p�Eq�N�r�!���9ܸi�մ�P9��BZ��!j8&o��|�jyoD�ނȭ|2	U@u�__">���Z�r���Ζ��o;�/]������W�xi0t��/X�V�b�$V�	6F&%��i,�6XI�)7�����\�L��V�&�J������]|M�B��X�֦��p�4��/�b�B�N~�G�&���W��p1|�����^߰���[~��,�;�"�0|��D��Gk�j�B�\W�t�WveK{^_�{U��S�ӆ��GwŮ��cn��#̛H������k��_*���R"s̻��e�2�Y����P�6��B��y�ߤ� ۬P]*��h%��`��'�)M)��|?��)��m��s}�q���t�����\B$Vb ��!�?����`+�YG,0ca5x���ދ�QBJ;$Z+Xe�E|1ֵ�jZU*�5����-0��2�{"�GԶ�g�x�N$q�匒���A�`�}���3��5Q3�`x�Ez���rQ�X���~ߚq;�:��on��1��<�S-i��}��˃�$����$�C`�8i�h,]�@�X��(�ׯ�bJ�^0�e�-�;�z��u?㡱����&�~g���Hz�kr޼�\�����H�d���:7�`�])�޵��>���;��n�v�ɕvxҐ�Y�+T��o���B;$��x�ʹr�Aaci`yZX[�F[6�� �Wd��D���R��H�����	�Nǟ������1m���G�3���阦�n78�JT�4{�c���4�l�tv�:7�"�p����e1���7�I��Be䯂؞��H�`
f���;{n�M�V~�9BtS�4#qSK���M��r���3c�P��xN��浽 ݶD�(c�����E�P�#NC�(�g��=�����x��� �dg?\��$���׬��9�lo
����
<��Cǭp�P�sm�i �������_7��Es�<!iP���My
��ڬT�20����=�
yR����Z�Zv�s����@w�.8� :�7��#J�-C=t�Y3U��lV��f{���l�@ ��\�=έ���6�C@�]o	K2!�g[A�����(fF�4�?��џb4�y��^�YҖ�ې�S��=�^��U�aPז��Kg:��J Głd+>ԥ���@��5v%�&��X�.�����|o�4w���UF�}�Y�f�Y��Bi�T���O�5���	��k,�ۚC����qy-[�ڨh��_4z����2����g2�Hי��k��˔(G�'�ay��`�'���a䃽S����u�#����-&`�E��Lf���9�������V���9��OeR�]-��\���P�ܠ'�x[&������Ȝ�vh�6ݒmv��E��;Xt�T�j�G����Yd��H�9Ťu`��OY������LlUQ*`F}�j�,6���dMRrL�c74�:Cg^���о�.M�3�׎vb��]�Į����B4:j�q�򀀤a�s��.C1�;)b�����x*I�TO|�V���'��@�-�s�X)~��������33��W�>`v&0m�J2�@���ri��e	M<v��u:gz'��D$ݓo��X��C1��v^B�y�&oF9��c�*�[�bL6b����3�I��K��j{�'�#}$x�����K���Yx�	=�����#/��:
c
���Ƃo��4|��� `���2����Ψ�s�W��X^���}`�ɴip�~k���޲u�P(X.z�Uc� �l.R8����T}`��Dϑ�G�Y|�;:�����������8���O�"j1~sC�S���B�2W�]��(yh�]Pq�n{��a�YV�Ğ�?)�YF#~Aŏh�\��Kp�r��>l^�V��&h��G�4�2C���W�Od���Ɓ�&�
��u���aX`m��i�H�Z��,���!}�u�#&_$	cF�x����`�>�P�@r ��X(?�fU=� +�4�m�i���D�4Ua�z��pB���M�	v�U*G�2��&QƗ7D[��\�������8gF{Y"�_|��������^�g㮐��T���Uc���e��菤>�]}��f��|��@R�����=Z���=%b��I�n��e�����R:����%��z�����Ċ��\m.PW�M1w�
�u�}J���\'Ka,S#���'0'��:��y6���E�M��c�ȏ��7�N*�X�E�Y�"��K��q��yUɅ�glf{rol�s̃��G3���QO�O'�Z��]���:�Y8��~.�n"���X������XA��?�iq��r���nX+��̈́���SS�
Bv��ɍ���+�������S���Џ�����!=6B��?qD��3�H��#Ԩ7�=eΣѨ0QM5u��}���m�vaN}.|j3��靕;Y�j��)��G�Ȗ�
��s|�? %C�j�2Y W4�5A�9��[�g�O�V��
�4�Sl�t��AEG���'G�B�"�Ł�1�7V����n~ѫo��R�}5��(^s)����bg�v�iQ��m�W����@5�ތt�_�k����d�K�xʸNI6(	!w�a,]�'�AaS���_��
n�l#��6�,�s�
)`WOط�!C�q��s���\���s"����8�v��7���x���H��:!�W,UY�;E���@�!��f¯��L9����K���E(,�������1�FU"[�͠7]kW9^�Jx�����5K�`B��qc�`'�^�U��_=��Q,�������
�t1�(����E_��^����Ծ��Ġ�nfEz�I<꟫!�а'���(�<do�:�@���'Xw�wQ`aE�LC��LJ����(omU��`�L�7������83��&��/˸V�K1��^k�dD��z�Z_�&%$��b!��q�"�V1���Lđyo���`�N)]Mk,�r���4�:���R��+U����^��[�yS�&��5^s����ZP/.��"؊{�����1L�8u@H��C�s�v�� ��������n�f���7�,+�Z��dO�.�1���=�֪m�DX��D�>=�P�V��3�
�ī4��C���ľ~2.��B�2���d��XÓ��m9\ͼ���8I��}��0��o���7�BJJ��?����� ѣ��B�G��
���Q�x-A�?��y�WK�Hc�՜��U��O�)���xo޴pXҥ�H�V��I[�4>�UsM6�ܳK�*$e(���m���9[���13�;� T����/kO��b�;���� �H#�{��%�]���L� �}��L�I���T�Q�b�G���Ob��3"�u(^R%��e"y��� 1�5���$%�:��G�C����\�eZ���<� ��#l��z��R��	�?a�F$�>�mI�C�ŦC
�6��%˿��J��yJm�$����L��qu��ýI�Z��4k,C:��\Կ�@����*�	��aw����/+��L�:Z{ZhV�ݘ��UgI:FO!Nz��H�����EM�Vn���,���w�u�O巘n^5�'Tzm���v~�M6=nŢ�	�f<?��}hr��%��O�Â�Ũ�M�,P$�Y0�'V��V���v,�N�F$ k~�)J�CKN��!N�V����t�֦ �Ǎ����A <WΕz�y���פ�f9ʛkuxK�B�L���慑R�RD���ͱ�>�i��3/����%�-p��
]�?
D�RZAɚ�'�ιb3�Rc�wU��ݓ���|'�9 ��r�~g�@� ���w��Q��@�"��i��A���V�]�0l���|]�?�&B�3��@��:bXk�p/2�'�� �w�z��i;�����=�o�-s�\����������-�ش���X�In�
:9�?h_&����4&c�A+�4��<\��r���$k6��(rʶ��v�k~Q�������`����ϮJH~��[�`fHr���Ud�m�W���d�h��uً~E�r���m���0�4S���X�4�6�p�s�5n]�:-=�&ΫOc��Ac��1Ԛ(��4��-Ht縺Ɛ�IV�Q�"}��F��9%f�m��O��:�����ٻ=śD�,#9�����UxK�I��T���`
���.��g�DH��0�r睝:xZ��Q}�� -��F"������p�>�ޟ�X���p�aZ�8 �UCqf�x.?����OŨ��3�x	Z����^��`��1"K�k�ZAѢ�$�B��>1-��wB�H�ZXv������z�ŚT�#�^��:��k��1������|�|�^� h;���V��EKt�p���|ݍ<3��  ��� �]'XB�H$��ґ���n�ڷ�.�j�4��_^�L�iLz���-į%�#��Ic��K�v	��tz�����n��J>�� 	��s���;:�o+ɤ�7�yj{�n`�E��PQ2����4���YQ˒j8���L*�է�P-�-�ր��J=�N�!{��)�oɜ�ck��S���4�#����06p�=�=Z!�aCv���ӭ����GO�F�A��4t�6��Y��?	U�%��4]X]iŲ��1p��e&C����c��Y1 .y�V�[�eݟ|�	�ݧ��_#�y��]A��B�^ðq��h�������[����U�ޏ�iK�
�5`��`������r�.������J�����L��+j�xK��ϊ
�S}�Pp?{&���P�˦%�`p4����T����6W�k8Y�J����|Oʽ�1���6�W�B���N�m�8��U���J��`�C�g��6x����kP� d�z	5n(�F���Uap�l�l;�ZϊE�#%��`�ރ�"*"����5�a����N^�#���}�*�:�E1�0`�gp����	�+��a��
y�Kf��=���3�B	+(Jb@Ǿhר�R3�h�8��fH���q��� bO_,u�z��!��X���T&��Pl;#�>�;����.3�B���ț�(gB'hvԍ��~�(�K0P�+H�������RN�iW�@���0��H;���%>p��76�1�����P��_^��lD<$���-�.�R�/��VɦC�	����+G� �[>��k��=��G4^�-�k����9ۆ��U+����M�ь�༜���6U�[;ɳ��e�v*iX,G�T��0��X4�h�������h�8�Q�NC�e|�Ӯ[m���ُr�ԫ�kdu.��ƿ>M���>%�.B�t9~^���?a�}�Hv�,�m��yPz�R��LrN��q���6l�7�ig���KF4`hn|3�Sb[;I�:AW��%���r��i�=kL`_�~�u�v *Wv���)��^#v9�%�2�B�ڲ-�=�mv�� �;p��ԙ]>�>lz��r�v`(
ܻQ��>�+�\�}��Dՠ��uoO��Q��,������rx �PH�`R!Q >Ij�p�0c�2J���s%J��
X�m��P��ɺ�¶�M1���O��R��O>�#�94�H~�ziv<�d����4�u�40�:3K�u�Ă��� �<�z��Δ͖�8���`�\��Q
���\@������NZ�<]u��Zx��4R��5�+'?�|�8���4ŏ��&'B8Wbk���U��mý�H͚��_�F�H�=�	!贌�2�Yy�Wk��m	6�����A���`�n�k�X�)68�	�ܷ��^d��m�5���O1�O��i�X�|�җ-���/fWR�c	�|�zCl��'D[`�������=��K��dM���6����~�jv�3_�ר�t�~��V�mg���\	�a���y��}����I�Cb`���<s��*���������� �i	h��T��а�6�Z��|W2dT/$t�n"�dj���j�j�@�|1��I	���`�m�kh�$+� �,eU6�Rǭ��=�|O:�,�q�V��c+w��6�CZ*P�-�'u��C�J9\��~j^.n�����ם��'�8�X�3�o�Z�R;f�E�g�ks�0P-dc��g�e�O����>S�&�o�t_V���.7�@H��Kۄ�I�-��@�]�����c�\�A^[�8)�/�R���~�\!����,aa���n3-T�EP�����E��_��릿�Fo�c�/ر4ҺWZf�Dzb�0�-��u
;�<y�w��.�����
؃n�I���6�wl仒�s�~��8����/�WV>�>p��u��
�����T���[��<����1�f��^�����sGT~�/�N�N�F��ȠSG���(HM����=��6�)���y��R'r��~r�g���t͗�oe�LV4"��ioG�[�>x�S�xOL��Z�-T!�^\=��I�A1���tv��R�(>}��_,8�&�V�ng8�OE�藲��2�ύP��A��P�PWHs��O*�͑,C�~c�y�w��\>�t����\TL���rc����Ʌ�Y��_z4`V4i��f���C��� ��ә��Я�!�T�K�g�)��~};��e�1D+@4���wM�Q5po�?O�<֦�?DS�[�).�+s��G,a�&��X����v���w��r)��N32|�:��:%zP{:�������XͶ.%}R�.��7��|q���~��RTWV�V�����}���L�U;H���������yy�J1��3u���w��=�ƫ^'��� ��G�
�_?c	>�
B�kgH�n��=u11_h8��E~pǝ�:�c'������X��t��a$���64qO���5<er9wg�KO^��/��J������Qm�+mÜ~�� �q6���׉5u�d�^����3J�ޘ��o�Z`�I�uv>E�X��31A��WM��fTe�p��O�3CP�ą�%<�h����?r�fq�T
&��b������͕���}�ɦ�_�஦�� W�|"o��Q4�q�H�(I���/�����%�)xt"�C��=a�]�o�u�qfN1O�w��xH�n�t,�1����Ŧ����"J�񬑧��L���.?{ʾ������P�{�E�=D����CP^n!��f:_5��.��L+8MP*�--��UW�uO�j�^/L�N:����N���˂��������{�C�_v"�Y���@0"T���n{Ŵ9/vJe=���<�M(2�|�k�M��l&��BD/���P.R�Z�3_�#�)f�@�{w�T{��z��2��1j��Y��l�b�1�ɚ2 �CY;���
�A帑<�'e �̱H�Ŏ�x�f�q�e)f�����~4�j�����1�E]<��=B���ʛ6����|�dP||D���0,����Z�d����/1S���K�~M�9O��.���mJ��ʀd�cAZ��H*&�������������2?�O���.ү9�@�S b���bd����|I�ӭzA���>��4n�@�7 �������� e���]Tm �<�n�4i:�� �lA��Vv:a&�j�-��]9�`�suģ�BU�EW
3���=L�G7���������i(Z�=��M�nH	0}��AOO��C�����K[}�J*�W~pd�ǌ���ۑ�(�+
t���4@�mq!����ω���r�n�$=ds���M�v����ka�� �;~��M#�	b�\�`��)�01��fJ�P�:�f���Lu������i��ߏ�0�779ݿ��A3#y�<g�O�v��2~�g7��Y�3�|#���x��ꬊY9�NP`Y'��U��L(I���T��:F�������)��:���UmfP8R<��a��}z��M��ۈ���~Z�-X�1�Q�\/���U��8KٗZ�����E�����=��N���<���+	�,VzA��y����`Đ�Ԧv=���j��;#J4h���y� �$I���C��-_|sm�g$����T��)����)W@���A�v�nR��Ѐַ
��K��mz���p�'�*Ц�v�E�_�)0"'�gg������<O"�(�����P6�q�e�q,Ⱦ`C���M+9�$j���7e��l���Ȕ�#4�5�k�:F�D���+�nbOg�X4Ċh�D�i꣡��҆�8��i[���,K',������)J��fq�"q9����{c�A-L9-CO�1-[N}�0���0t���=�6�*��cd�2_\O"�>���6_����������1;Z��:㧄e�W�\�%6S���_aA@�һ�4��>G�T��Kp���逛������vע���VT�����h1�hѲ˷���*�{6Wb�#�;K�����6�W�B��w�	�Y4�����0�Xͥ�yn�@�������J�9�;�������_;���(�w�rϣ���|g�(5_��d��^GNّrh�5^��$��G�2?7ӕ$g�Y���:�b\G�)J�k���|��fD���NA-'���jCw�+�rZ����i��8��m��4m΀��30U]'ZX�ٙ��ǵ&��j���V���R$�e��k��� Q�801�v!��|eyѵ�Yep3V���~��j?k�7F�
�ɔ-�P51|.r���KV'�c�3SW-���(�uf��3~�gM�ǲ�:^%p��T~��G7�Ł�\v�r��O~k��t��#5[Bxh)g�*b.a�U��Rb?���s�h��[&ņ'(B�Q E�^������F""A�:uv�h�s�V5�2�ֺS������P�f~ߠ���z��}
m�����Y������{�le�+��*n����ﯗ��*eh��G�6=���|�z������s�-�՚�b��:��)����O�]�~'�P�:��[0
%|�٢%�:�իq��n�|S��{K�O�"u���bg�EP&�d��1�t�q�fg���Z�N�N�6@u�H(�/���V�y/�%�-�4��F	h�1s}��_,�.
$Hc��@	����+������_u�J���	$q ��R���^ �oo���rJ�=���ND#ؑ ���TOD�R�\����X�M5�2�tJ�Z�Z���PB��qÐ�ޜ��ޱ@ݐ��j�ؑ�7?�7.�,�C6�V��Z�)�GF����N�`����?��8֖	�	�1;�P������i�����Ό�}��'�~_|�L/q�;1�����^�s��M2���E(-���^�Y�"���5��y��6�t�1�8�i[��m\ȳ|�N�r���[�����0���5Q������my]��U��s����zu�� ���ȑ�5w�[U.V��7�Q%ecF�d-z�L�4ס��ACD�.A��o!8T<fm����˅^��]�����\r�����>6k�a�aM�rو!O+�6�%*�֑x�0B�0��߆��M<���S8ێ:�U����v?��3%ʺxb���Ό�f�3�-��;\ZO��'�3��;�lL����'A�Rn������|>1b�^�L	��i�a��X��S���H��m��}��_J�D�PO�[�@+�r,�G�xE���"ZQk:C�{I5�~��������(±1E��C�hX���\M�8��2�!R�LsA���ڍ�*[��u�4W>�[_�`?Д�)Y��݊m��$�&yҬ-X��5y6T���K�5��G�[�����r������}�J����_���HQ�ܵj z��Hy߉�}���f��.}/�Y=5��� �,o�bz8���o����J�ם�Uة�׹{.	�+ݏ��������T'��@ʳ��a.�;�s�os��Ev�U �	:\ y&-;a���R�6�ִW(�+�9��ae*k׆���~��遛�6k�r=1U*:��&�@]g
ym���v}^�feY.��$\��+fT�5�4��0����P� u�,f`x����W�h���j�aK:r	S�p�uu�;�#��Kz";4���������*�I��>�Cg�B�7="�Z��lF=d�&+yC<��o}b+��!\����As��'Ѝ����2�G�_���]�uL[��	���f���\����@�YR�z���^%[-��M�W��E �,�O��J�R�V��Jgv����t%#��(:9J�����zq�m���V��h��4��]��DS��*�I�Js�a>���ϣ/���$���f����MD`1��]��j$�T�������D�I��c_�8�c�T��>��,�r�Y�d1]Pa��"�[�8��f[���~�[��fC�%̭�ɶ�$�J;"#��Nw�/��%\�g����N�,���א��u �'ma�w4(W<�_�۝+����0l��j|��7\��n/��c@->��2e���.@��;���'�J50ܷ����V�,ى�bQ�ղ"���1�U.9H��/�WK��nj�ũ0�d��q98�G�_�����������+�"��v�h[�o��TC��Ĭ�Us�Y7#��#�RM;bIt�27*_��f�D�H�"�q���[,���m_Bo؇�ބJ��BQ�	ߤ��<���XXƀ�oݢ�E&�$�[��Ъ٪��#|��[�������[�l&:6���U���bYפ�Fba�7�ܱҧ���-d�1zI�&�}�#�lX�4�ZzA��Z>"ʉj���"��z��,�w%������*�s	Z_f�Ճ2��p���To���7���Ih&`��w���՛��D��*����5
����:�X�W���@{�G���:���gu�.�AB��X�b�$��������Hʗ��$)�	��t��Ո�J�nr���ަ06S^�W�}J�*g��_�R�8d�R�6�5��j?C簩�Վ�-�mF��G������BS�9���Y�+��^�rzg�Sn]��Jm��5ѓi�ā*emH��%��9�g�0ME�7�
*{Sѐ��E����:�yl��J�Y�-'���OI��z ��L��7���Ы�XɌ�жP�q�P��!�;�xd����W|Ю5PrҚ�{׎s�a��:���3�0X���o��K�-�N���c�_%�`�2Mb���[���"d���#"�?';�B�����R��p�&f��J�򞪔��qЈEь0H}Pm���d������k����Z�GK�'�o����LZf�[��ſs�t'�����SF�v�j,4���B]T,�����ե:�4-�Y�$�O3a�ޖ2;��(1�����qǷԱ%���9�+8"��A�����%��uD��n7�p��sW�\���h&��a?��
�N���J�R9Y��5�D,hI_����s�.�!|PR�PML������8�U�Nx ����I�z���d.�DK��������*D���U򱵈a�C��5��N=�� T*���;�ˎ��b��S������@��1�p��Z��	^J�4q����`�3�V�]p���Ͼ�|;�s}�_�H@���
ۍl�,��R����If+o�Y�=��I�������+��rn��E'4a�b�9B}�,��w�z4-٧:�;Щ�nZ4��7.��]��4�h�����������V-[8p�ɒz���"̒��UR+^)2?�!�e���?���3��*6��!�d���~	L#}��D|-E�\=��HZ�Ih>j��=��i��c�l)r���]��n;��#Kw��&�L숏��˄Ƀ �F-������'j;�-8���ێ��a�?%Ę��!(�.l������B��b?��^�Cc�X �;�9Pozi��,����)h ��ܼ��?4�ϯ�l�bm�3�+�dxwV�����H�&8��(� ��2 �_�!�n9ӂ&��hXF{3��8�Yz�zV�曁ܵ �H�:���<=��7�d���.�m���}�8����~�2�	c2@��|�<�_�����.�Kp�����Q�Ud��B�S73������m���vE�oX���U�ɛ֫��ÑR�� mL�iK�ls�cI��;"�.� VB�Z���s��8���"v�
 ��,� *�s[�c5�,}\�5��~ci��s����K@��E�A��������*[�R��zSP��DU�[ef���p��F=��^�Rx3�I|���˝��Ba_�(��t]ν�V�dg���c��G��;3�4����z�����>p�Z=L�`&���!��-�g�O,b�۵��2�����6��٧}t *ԡ	��T���п�g���=j�ϒ��:�8�?Ύ�حh1��,�mZ����=���<�Rb,�a���-2��~%�z6Mb�4�(����$�/�����q
�"l �N�U�h�ʚ�YP9p����\�;"�c�;x���w�qw���C�"Q�H��ڔl{AT�z����\,�69�J����Ǡ���!aeh�Y0h�떪 ��䰾
5f�,)`%�>D�݋Q�
�=�#>ģ���^��Ϋ�íZ��D5�2+���#�;���߁��y��d���������;��\xނ2���^�E,�0,??
%�:��L3ퟲ+vDK ��B�m2�I[!�J�舅C ��U��HŅTºy��av�[��2�ݪ�I�>u��N~�*�?��������U�'.�|�>���+M,�G�Β�HO��	���}�10f����"� w��b?eG#�cW����钡�ku�q'�tr��[f���@nH~�4��nwx0�ϋ�VSﾷ
��	��Bnű�ll�[�q`������l����Ʈ�o��{j�*�$��.}&$�٫�vy�}�?�;A�*��`�sL_�˯��V_��3�L��N9��ȋ����G�\{���C@j�K����e�$Jn���Z� ���F��$$zP��*��J���n�dس%�ۋp��fGU�(��`�o����Q�t�Ħ��
 F��q7V�	Nbe�¾Ǉ$Y��^/U\(m�5���W-�^��A���F~E��P���Z
o>lb� 12�h�����WY��H���2f���2��3(es�������Z��>B#�t����D)�Fa�;OJ�7'XR��&�O�c����NG��:����������#Ees�0�ӿ5&ˤ�?POX.�o��	��yQ<�,!YAR�}�L���b"��q"�1z�*  S.�S�t�;M����i#Ax oԊE�����~�ÌE��ǿw������|�O��ؙ}�K��笕y�JM�x��j�Rb�0����<s�P�A��/k�eX��wZ#�����d	��8k�|E���E���o�
K�^�F�^.gKh�c�_�6y���6����%ປX�s����?������6�O"���<��7�_�x�Z�־��(E�O�6ޜV���J;	���ܵ��Pʞ�j�����g�ht�X[ߞ���Any�O�vv�jw�'�7m�u�=u����Cte�>���"�)��-0��jj�F���3p@pQ�V�"����i �,4����_�Z�U-�@s�Y1$t4�!���ӷ��ɴ�_4�f�N=���âw�J�h�	֕f��u�׻G��@�В'�Cq��c4�gS9D�A�������1?��/Z|L�S��d��������hGd5�����:x�2��q�,����l��RD<nz7g��T+b����v@��$RL��:%��"޺
��Xɂ���+��3VYL���$�(�=����ݸ�᳽�/[X���j��I�T�,w�ti�8�j��|��=���h�c5�Ad���R�U���b�R�3K���qN��^Y�?��跳XxS1�p:�ӲLD%��
�ÿT��J�al~�2T#c������ҙ���R�O�!\H�LU�DeJ�w�yQ<�K@��ʦ��_^F���P�3�SI����6�(�}3�����-���3�ϟ_��4��)�����[e��:�ƺ�����UĐ���-�Q�M.�����%?D)E�N��뀵��P%��C������({�5�T^b Q�\���q3�@3il$��}+�(2���L�#�AQ <�U��8*A��(w�gn0��77�R���Y���:ʇ�CC����#�m�r����s� +5Y͛^K���`�>�s�U\<��^�3M%�?{f��c����b���%�
�.;|�9eY��VJ%X��^��H�ܩd��'i��2Du���16v���\���@*�;C�W9»c��H8��"Q������/�g�(�ls�Q3������x)���9�))��2@�5	s:�*D�_�C��<P��o	�F�L
�;�O@Y;��:���^�J#�%ìN��ȃF��i�R��1M(���u�Ӝy�[��4X��<٫|�"&q.&���I_�"	�l����9I.������K*����0pkq���]Y���p�ki=\^1���*{��K	.�a�d�st�c ����w��'��N�_���gec�M��y&�kJ��0��n�F�}�%�q��V�aN�����Z�ܪ���o���.9���_@ѹB�����~�4M9��w��_ J V��8V������+�Ϸ[e�)vfn������;-"�/t]I����~�>d�e�gmLd�fG^`6�%k�# ��<7^Ю|�A�'�̐���֞�{�$�D�fc��� �v��-O�����*�/��Yw=@�d�˻�%3�~FD���.m�] P�w���ˏ�����W�� 8y��N�K��h��U�e3a�?k�C$���2)�S�m��i�衇.8����6�ͼ�˯�C-"QF~o2�ہ����52T��)!!���'��O��dU����	wK]�
�v*N����f+�I`��������4�&�1$ ����F�rl�s۰�d�p-�Vao^���(�geYI)]�{�Z`��"V��ry�7��1��;�J򑁋�*��?�ԂG�\��ޢ�b�P���U�L����d"�P��pР���h�I8��or�.���L*��mtd%��ۊ�}�i9 �)��l�K(�7��"�HA��Gr����f��RQ����K�䇹?0��x�����O���2����u �����LC�(�Ym-<�(W?�[�5�ȯɢ�	��gL�{k�"��(���.�|�`������L3�v�i�"��[���IS��[4ٰT�Q"Hsk���'���gKB�F��9,�+�{�����B���0܈�����j��LY�J�x�X%��g�����W͓�׾�@��Bզ���I����֣�	�\.ZK�l����5���àm���#��O�Sά<M�;c�lV��Uc�Cz�;M����EX۶po�3��7�'�W����ʰW�9qՠ��xu�|�K��8�Y��/��8n%_w�/�Q=�,H��x���5�7�{�yE�U^m��~ȟ��oZ�V��?hTq�"0�'M�S,��-H�A��e/:�&�urj����jR;�psyM��j�2jwciE��.ȕC?BN�aձ��(�^85u�q��Ӈ�YX<cK���T��'m��:���b�7���4B���7=�^���ɽUδI���7;�: j<���kġ��Ժ������H�����/}h�8a��+Zƃ���S��Mo����6�3���{�7��vhTQ�9�A�D��V�F�#�wՑ�����O��@Xa���o�=��i�D�[4/����w
���(���h�$Zxj?ҽR;[<�w��7A>�R����\�wdl��Q(h������\�"
7K�U�#��ʌ s�B���❁i�~y/���m:�����؍,�����S�e���k1�7v5�Qɕ��+���)�����T��őQ�>����7g�$���e�VB�3I+�N�k��\�Y�>�J�@?d���9��E�W�{ ��af���} �����!a����~P���|���V*���K���0�c|]��FT!���xhʑ�ۣ4��:'W�o	�h�j���e-��'c����R
���W�e���]v�����������c�J����)�&�wB����NX��Z�$sT�-�EE���n%ͥ#���^a�@�\��3�� rP�tp$�����*)0��ETw���`lەEJ�-�`���;�򞍒-���m�Y�O|�jW��ޤ��������|8ƻ��(k���g� !�@�%�m	Fݜ�I�o(�0Ȩp:��Ca�QB��m��㼆Ⴡ.$<y@: "�3���*H�
%w�a賏_�9��Y�ÄI ;æH�L��(����O�or�95��
+�_�[�"`
�8����y�C�i���:QeP�<n-�x�5a�BH��a�4�PĨlʫ�S��?�<2p�9]�pCǹ�HߛSO3�Y����@L��G��4�'s�x&%.f5��;.Z_4b��o�$��6���&�1f�z�Z/��H	g��YL<h0kJk���}Y����+F����4�;`�h+���&ѐ%�h8�UH�ܧ]l�.תv�XU}m#�ݖ�;�σ2�:p�����6r������ᇄ���x��m�@�%W�9k����2���ҧ�M���{�l��lh?�sp1�2@]�/&��p�f3_Ջ���4],N���<l�뜠���Z��S52)�E�S�fo�"w�&,5tw��(hhp'��}��[�
��v_ܯr����J�y��~��5�Ċ�g�[�ը&U�>��]-�}B�+�G�� ���Uʳ3�D��RN�w�$TT��L����}�t����e�J����)�ʛӢ�	�Ν��:�^�����K�=u�����CW�#�ej�*{�&��k� &�����Efk�=����E�2�h�̣�;�p~h-"��aƩfN�������[tά�M|`�9>9닰�K.z�Y�Z�t2kKwM����6.����=RY�v�H��Bw=�c�d�����=I;n�*6��|y���!�Su~�-��86��>"��<������W�z��?�;�d6�+���K�%N�Z��O����ہ6���������9x��y�OA��r�,� psF��W��X�]��B1!�P�wQ�K�G��ޜOS?�J��d!�b?�-�tQ�ǔ��)]ף�H$���ﾏp#=����O7�,58�g �����+�U��,&zs��/��L�p&��	b^���=9��� ���H�3B�"&��Ev�o�f@�q�^��}�:�j��w�T!ô�I�T�ֹ1k�UwMB1��0K�>^ac��ʦoj�` o�t�����g���[S�f��]��<S�AQ
;O�U�E}juZ�7I��i䎪� ��,z,)����܋�P��>[�ߒ�[�߱�۶7�;�B�,i^� �bb��a�u�	}��X��D ���u[#��P�x�fĚO,�7��V�
&q�0���@x�df���x/�C�&��I����ϨB�u�g]"ϧ������}XK*I��z'B��v��ܑ�	�H���A�����#,S�Q���L�
Ë�J��\=�}'�*����(��-:�a��(�[�����"zReH��q�-�\3��/�Ͻ=�mv��x���:{;��#����;���RU�r ��
�Sk�-4,.y��a�ۓ#sP~�V]8�9����7���{,�ڈ$�n�O�"���Fu�[��눂>:p�Kc����(:���mo�Ų��[����#N@vu,�J���GmՌ[�4���e�����K�o���&��ur���:�D��Ҋ_�[��V"J����U��I�y�GB�?�;3�&M%9Q/�L^Ͷ����U��c1�1^��z)�Y��#u\�+L��� ��E�ہ_�����IwG�w�7�O�R6)��ؓ����j�T�? �������[���kF*^�-�#y��O��87���M�vw5��K�3����sta��LyD��:���+���M �,�	/a�(�(�prR�'$�U^���� ��rz3�����Z�����n��G#�|
�����zS�+�:�3�ؿs���� [�7�>X-i#t���-��z�M�=n$"s��ß1ǋ���FEXG<�+�2���Ug��\X�����{=ڰ?1w��v�xQ�-������a���
K�a�ߤ6���y��g�>��[SC��MKHzǚ�����ߞk�$�bo�
�w��P9�y+(�7��}w�+F�D�n������P����A�� �HCV��?A_e�t9�`\���SH{�F[}L��{�Ɂ��+ubg�Ƀ���g�=\����,���詹�D`a����b�O{���ݚO��`I~��X�w����-�+�Q��q�N_p�z�ޒ�� g�5����-g��z ���ۜ��	�s��3��h�>�1v�1�
���Em�gTT!>���Y#۔�T�RZ�V�������|��'ͪ;7T�ꨥ��r�"��ј氿��ZO��ίQOi�O!^bx�q�q��Ҭ,׾:�$	226Mv��!�bt�g�A<_0��|��/���Y��o���S3hX&/�&�X�,i�tt����U�#�t�-��w��c$�#�KN����0�dL��J_�Uw��
?�G�a�irD��6O�pp�-����"�˙��c��3�(�V���a�~o���:x��1��{"�E.lwW�z�b�����pCrHh�h��,<�����Q�`�E}="m�HסZZ��OD�L.�;��%[��WY w-|��+���d�3�O?]��q&�;,J�%a)�Z䘇zH*��1��*"0Vio��=��;[P4q��؉��@J;2˲�{&��O���%�9?'p+hAdSq�n�����-�����i���@�=m�Ӟgq��0,=Ğ �s ��z�?M42M�9�]2��tI��gb!p���î�YG�*	`>�Mɭzo�Xu�������Z����!F�1��ɯCt*`Y3 ��b0���r��OY��=m̾�=p��w����@ި�)+�|:���H̳ʏQ��x�9��x|�����:Ψ��"9Q�u�_�������xȣ��h�^���"�+Ι��C��Y�J���:]�S���D��V'h�4n[�A$歇�=H���X�Y��5'~aCh���MJ?�C]��%!���9'��吅FQQ�N������o༎sf�rδ��;���7(233��`b8=z�@���>�a͂��(݇E��:A�gP�y
Ҝ.Ѳ]jF�v�x���J�J~4B���G����#v�-:&%@���U�����2D<�;-�(^��x�g�$<��}�o�z�c��5&��X�"Q��w�AL��-k��eR|R��l��K�q�8G���>��-�.�����2F�����/�6&�XY�	�%�%E@��P���^�T��+�O��-8� �tM8/�K��{�ϳI{���8j<�mG&N!p���������|�q����<�/O�����KZ+��`3����	���IM�yޝ��Y��;:s�/�9x6�9L�ͦ~�+_Q=X��%IPv�DP�S��P͹ZU>}�!����J���&@���S����XZ3�m�+�W�x��M���$�?�G\1�Y�哯w�Ŷ'���@��~!c�Ɠ23�v�:��/��[Wq�^<�t�~���F;a����Q�;��ڛΚ�D��C�͞]j_ɜ�����H�̷�܂�JZ{O:�Q�X�������̣���٦.�y��Z��5]���(�uQ_�T6��!���<�����,I��pVݜ����iaB"37�3R�U�T��t;�=��>>L[�?��!/������D�w�y��B����a�Xq����?t�������77oevɯ,������vDx�7r!�,�W"����R𘯭r����C���ae�D
�2ǪKC$WW��	E�upӋN���?;�<@q���F��m�~��T�=�X^I@�����/w�mJ�j�;^>x[ :���D������%����'��QA���dn�@��<R��������=��a.˩Qzo0��rʱ��KǍ��Ƶݻ�{�՝������`�1(�&�fn%Kq��=���dnE�$!*s5?�Rl�`��S�32'Q�z�y�p65T�7H�V��Ƒ�ܷ�Aտ�,����u�����[��)��?�4�w���臘d33�vU�S'4L��(�o�Щ�w��� #ov�a�S)�I@0�a?��O\��_��sWÊ�F�+�~��;��A$������ub�M��_�<:�?�y^��.v�Rd��`��-Iq�a-��޿�T�L��15OiF}�/s[ ���3h�>`-��5'ؔi��׭�	�ciN�����|�թ$~���R%!&ᐎ�7�!��B���W��Q�+�#м㇄ }��G��$\4!R�{3��R-Q����
�ٻ��,��)&5��|��-�l����:�d!#��ze��`�4��N�D*!��9Ln�6T��2C��q��8���б/L�MI@�A�����.�2>�p�V��n���U���V�!��˫~��6c#B�l3<�#V�`�p��h~P���2�J:~O����`=��Ε��n^3'�u��i/�)��9*XF�Tߓ�AO����O�=@s)�ޘN�Nj���&�C��N6_H���d"��iM��F�Ы��aWS��\���2�Fk��m:Cϳ{�&'��w�Zb�1=	D�0A��[1ͽ�q��E�T�O/���O�ܼ�az�>���4��1xh���P�.�{tѽU������@�(���b�����?��Q�����Z}u�)=���y�KR� �K��P�f蓚��id�Ak��F��N�dS	hG��)������iՌ�����d=4���LXq�<�fĞ`ig���v�����e����ME�q��G�T�yc�k��G�_��� 4T�V �ԣ���
A� �����؞��,*	/E�׏�Sc6�#���[�lU��d!��G��"j��M�G�B��7�����|P�p���.܉ �`n�d���}Jk�N��F��`�$g����|0C�6���}�R	�j�:�uw��>,�F�77��-��Z�R9�;�&"�і�p���Q8�7�[{DӘ��O�H���v�"� �؞=�aܸ�
��hxw�����G���^���C��)�xE,D�	)Ç�**��7L_V��H����Slp�p��|�aom�J'k�tmMyxG���U�X�.ϋ%�;p�D&	�5���b�BY��;���젝��]²���$�"�Ĕ�7��cD�0/4�l3�����ܶ�*�Q�0�f#/�#jfH26s:�<��r�����T
�N<)i�nwyn�7-���F�BX��I�?/d�:0��_!��bby xX"��։��Pݬ�JHv`uT(�u��Lه-���~i,v(;�ut��4Ǜ���5v��'�$ї�����^��X��6���+]�ç�G���.J�T���3��`��^�x��5��X4�u�@Q28�B�dey��pΖ������
����sST�n��s,*f�,Y�5�j�� �:�Zw���H,�򫨎ZS�|2�^��^.ɾ9,b?��R����=Ev����ʹ��(H4�yn��3�d��v]���>?趏7R�IV����B�1��vj3f�T'�J@גN��VʖiV�\������Ryè����y�h����ou�b���Ѣ�	6�\˄�����h�΃��� .)kl�?�_Ya�
]r�޾>2@��l1�b����x���C=���|�o$d$S!��hm։ �C����̉�!��*)��s��{��$��ͻ�N�*ӄq[�(�ZM&���<>`ޘ�<�p�Č��OO�~���(�eJ�;\d{���n�lC�h�AfEr�Fz�\G �@�P��_`!@I<dEi��[�t ������B}�M���шR�)�2�hO,_��9?J�&�S��m��GD����M�PX��o�ɡ?��J�qߎ-���r%�df�L�gB�x�3*7�����,�&�?�O(��N�(�Z�"���V`����ЁA�#Oà����_zl@�jL!�A"\������i4**0�Cvu���툿�j��{J ����nĂ�����GǹB?�;Kx��^F`C�X!*}x4��k�ཎ�e8�;^�G��n�0T��AJ?�ݓ�m�:"y�o)�EH�T�y�m�<�b���	��Q�֭@�n'�9�}�������q���Z�ω��DN�M��+S�V �$���MY�9��x~-L4��́L��8��e��14
z/KB�*�\R�89���a�bb��em�9qN7>���-Ls�ݕR{ݕ#*�fב%I���\�u��;�Q7!f��gkU}�L8ވuQO.�_�h�)=���(1X�R�Ne	IN���}��g�~H�e�#���B�SKY��!�����Z�ˉ��x4�{}kT�ޔ�f	��%h�]�n��9���������z_�����7	�y�����^Q���&�Qwy��wG0r��ꨩ�0ta��I.�[9�����Ε9�����x��n��j��%�t�����	>�^���-����:�r'�"��W�L�=����b�6�z俙�ٿV��k�E�Kf#Suسdx�����,��U^�TC������N��q������f[k����Y$��.���9 �n�y��� U9�<��'C+T�����y��,z���vcE�FHfx&�TTE�x��Ks>������LxC��Q"D�W`�>���/�P���,��Jx�i�p���+v��eELoꐃ�Ȗ�M}J��?����CST���Č��:ڿ��i>:�LVR����?��5zb��ӢN֮Q�!ͨt7* ��ޅ���J��
�}Pv��@����)��BE�����lL(�٨�ʁ֬��f(��2��aw�
ySjq'~L���5d��.V#Q��gɚ:���lS����6������،׏)|���������ܯ�l͂}jX̔��� H@?;�j�K.,\Y���\X���Z(O��z� )�P��߳{����ې�c�s,�3l	��X
�տN$��_�?X��ؑ8��]`���;@\c��ac��������W�
�`��3y���x�&`��#\��9?=A���5.�$\|��4
�>�X���Xyݡ�[J�)>{��ɑ$FIaP���%�c��⫤�����o��O��֨�7H��{�\	�	�g<�4&e��&��W�&s�
�7&<msIW���T�=K�@�m��&�~��pma*s*�q�~�O�|���˿	�,��}}�n`�A����/�w3����*}ɳ�G�O�ܾ>3�C�&����-����I�g����ʷ��ũ��� i`k�:Uj����&�sS�W������Ꭴ�ۨ�-��S�Jx�� ���<�x;Zw�ʩi�TǱ���1p{g+�K�HI#G)�u��Гw��r " I�O��<7�4�(�2O�C�|�F�2��YoA�2�TZ�SFϑ��Db�����Y}'�n��wD_�֔�.�¨�{�͏�e�����Ϲ��Um/ӻ&������=��ѾId	��������C\C�Hsπ��Au3�}28���B��B�A=ڞ��b���;���c�V�)D�E�z}}ۈ�&2ԝ.;)�dW������ظ�m�%Y:�+<����i[�jw�0^��?yN�'w��V�QM��kO�� TYe�Z��Ζ$RC�1y��n.(�x��M�#�������C`Ɂ�\�!��p�TA�>m��ͼn_1\��⾢<�S��Kß�eF���Z�6C_I�X5�h~n6�R* ��%*�=F�)�%���� ���)W���(3�kwI<\?V�TF]����[�8���$7�6=�u��qa���>�@h��mLtG�bVf�3�P�l������~T=�]�W��}Õ�7*s�-ް��i�̙���T����#��;����I�n;�sP\8M"���d�}����BSНpm��]z�'bQL�-6t�T�q�̋�)���r�^�(�(
��th����4e!(����L�c&������f�9u��{���R���Ӵ��н��fw�W�3�� ����XP	�:�z���5`9w��K�G����Dɉ���΀�~������9\���<-��W"�i*��Q�,�,�*<"��m2P�$����Ҡ��Ů�Ee%}�Ȟ����{�g}����繼eC��rGZ��V����J�-���31��\�nq7������vn���:���/Bu��Հ��
�)j]����>h' �JzVD(�Ʈ���!���4Q�i%*&��n�Iq>>�0��i��l0%�kH�{��!W�)���-:��bˢ��p�^�6��j��P�����l �eS3~bc�7v�����|�\���웁pw�m��_������8t����k��H��������<c_4��w��HR�7�8��GJ���ZV�Y����C޴=�P���FN��1�|^`׬>�-�hL�>��?dD,� W��U�D��,��D'���4i�v.����Vq��њN�U��Q��)Lٺ:����R/��&6M���<�$�oi��+��r<=B��[��2��nz�Xi�g��e��P�F�N����o���=��0>��Q���8q��E�0�����3��̢l}K}�EZ�3���uQ��qֻ��u˭!8�Tl@?Ch�/$�+�ǲ+�X��%,�o*�;���*(�mXB��4G����ki�t�<��0�E�j��Gb3�΄�& Q]�����o�����-uw�Hő���I`�Q��|�4��ބ2�aV���������3��1�N`�I�\5S���-���5�j�x��T>���}|�-v�fW>R��?�q�0D�
r�c��]�d��w��Tq�v��k0��f�#1A,`7� /�a|���/���^���Y=�B� ��$�U���N�LIV��"��\� ٲѝ�a�8��������.#���P���f�oH'��� :ը������FWQ��1��DT+u�PYEuG��h�-Z��,P�u������H���8S�������0>&�U6���ڃ1�*�ʂ���� +��#��B�,�̉͠� mQ|'���xdP���J]�m�r�gV>�Pn�z�	W0,p��r��?�m��K����:�6FW~�A��z`CDy�#�!�";��⧼J��w-�q��U9��y���I��X���g�N��i������F�6�˴�� T2e � �
`D�9�1�+��A��t n$�����Ra3e�D��esa�w�u����[�h��c��]#���z�]�T����$�{k� ߁�7 �>褨�Cg�(�v��5&ƃV�Z��c�V��)]<*�eJ�h�a�U�Y��0����Rm/ ?�$:�1Ą������p�^$��>��4$��fC���	�r�瞻�c�/d�I� ���S�D�x�`�^��#<��4�=q�<��g��XO�`�Ǩ�P��]&��x(�h��4�o��ٸ���+���mңІ}K&Ǝ�ۈ���ff8�P��v�i����w�{�m}�A���͇V�IF�ه��
&�\����:DK.t'3��p�J�B��;t}���m��+�K*�͔S��s�)��p�Q/�e=���*���|fsI�����Y���.���}�%�#e	$�� ���n���k-OyQ��#=�z�W�<8޵h�)�Ӟ�+�U��H����U٫I3j|�^̴������,
�nQ���$��kq�a�j%O���C�7G�:�O'���e�rCp;�NH�46M"��
Ĥ���������8��ɉ�k�`=S�?����"��<�C��T�?��6%(s��Gq��WN���� �3T��r�N���>Ɂ�[���o
T [�N�:Ң��PT�dq\���`ݥ�3�[��J��&��;.��9�G���x��ݕ�'tp��C�����{�pca[O% H]s�
��Q�S���8��XS��A�?c�2���
MI���J�Ww���	�n)��p^��"�l������,p�7�����ܟ4��_\���S�1_�=��3�;��oϵ��Ur�$Q��T6���?���!u �R�����&l�R,_L�;�*�.�#��L\v#	���d����)ֻ&�D`��%��yP�N�F;b_l���Y=�sJ�/Ԛ�(piL�H|�
���_�0�M��| T"��G��#�������AL�Ts�U�TT�^	�l�[�?_��6�������a[Bf:y�z��r�9EJ":���s94�?;��˾�{5�B���ZG])��Y��@��P��ׂoL�?���?�~U���bm^?l��Gq$������hEl���;�o%��8Z�{��k�4$x~�A����HL��D�ea�%�aq�-�8oXi��4~�^S��ML�Z#�|}�tG�CI�x�ԏ� /d}�ǖ9����\�&�V��S_�"��J.��8Ʋ���2}�|�0V>�+D���L�Y����r�_zmҼ6��Jk��q�� �a�V�h��c�(�X�M/��Tp�O9[&���$�o�7'z��Z^FUG�xC�`#��P>��r�N�����;�����w��ƙ�
י�>D)��C}���������e���œ�A��xl������WZI��hXon�@c�H`�z�V7%eSco��}��@�d�o�P��`<���j�n8Զ^�#�c�AM��I��j��l~j�ɟ:��֞p�5��)�t�C}A�⢎z�^�u��iq��<P?�>��b�����BQ[^֐�}F���Xm�K�w���x�k��l���(�i��##�{i����O�iW5������+p�����}�-Z�;��+�po��ƛ/��C�9J�(!Ǩ��y0����qxƄ���E���5`k���BZ�m��QT�x�s�yT��n�W�p�TFɧ~��<g<��S����� �<�&Iw6���X�鹳 C�"�e��L6{��^��WGl з�������D����iF����/�И�bxEڋfI�_�7
$� *a���p�C��2޸�J���0��D�]�V}�G�������*�]�$%���8�Y4�ST��4�j�S�uc`�B��+��3��
�z�;/K��(�bY�m��(��S�H�h�אIo�
� VZ\)�{5�4�������-@1�X�*F�,��!�Z���n3,�5@Ҷ�τWn%� K~�R�ae�m�0U�6��a�K �|Q�Ept�m6&��9���7}��'1��~[l��r*��21�sL���Sgg�ĳ�HCd�!�"FK��3ꑋ��!E���CӋU�iɲ⌇PY��(��eo�S����WX^��
���#��d��D�z�̯<t�����ͯ�cY%� /&�W��UIHq�'�WB�ʂ̬����2ڶNIMZ�ѲX��}����e>,�Ec���@�!|N!�W��0"5��U�`��nj�\0�Ga8�w�׵R��ϣ'�0q�>Veq�C&���Կ�L�}�=	�x}}�@p�}SG�vH�sT?���&����ӉX�jl���*��Y	�#g&ȡ(5���0}Q��M{dbQ"�Ӹ�g�{����<�&l���7Hr��\7�I�j��T2+޷�������v����>}��acBW����oQ5��j�f5`�GҴSݟlU-u��W�I`.�����P�c�9��y��&��L�&Ǯ���֣��7��]U��tV_���-�x>��/���H2��M`�o8�QͲ�~�_{S'[���D9�!�i��.�p�[QS�M~�Q���߻)�.�~V�#�4Sz��G
\��#�{Y�G'c�<�n�uA�����E���=������B+�Ľ!�"'��I!;~�����_��F�� :��4,Py\|���X�m�� P�h�o�-���g�M�*�&�:�ж���Ahx�j:�"8�3�R9jek��0.>������*�Ԗ�M�v";�h�xO~�I���% ��3Wb+�(�ܷ���"/|F<+��bY4ֿⶽU�F�}���s鑚W&n�g��J�͂��'3i��*�� ������/1�L�c��Ԗ3jZ-9{X:�U�� �#6hus�E�x��E�*�,.	�<�Da��IN6 {�汜�p�.{�
R��Wn|�0ӎ���������?���0���o���	��$n_A����$�
�;mS����-|U5�?��'+�2���
!=�z��b#���#���%p�.V�aP$�ur|�l�'���x�^�֓�H?S$�f��V������W�y�_��q����>����|-K./܍��;|d�w^D��BQ"�[�|t���y�w�����޾�/sĆu#^��zS���0�4�Tw�Ѻ&�-�%��=�l��2�������R9݀�%���,n�����z	�BrmX#�Աk~�\�i��+�[��"�$'�y!���]lգ����H&EE�\T�L����/�=���l�`g�<>�������7��?�zʛ��� y�.�Et#�0�g\�F�ա{@h�9�D�Jh���X �HBz�L���� D�7��]n��N�qy���y�,B�ͧӖ�&.
�;��cc+����X-h�+J��5[
��k��Z't��zQV�PG*�����$��葬��|��)�#ۨy����P�D������H��@�^;0]+-�X�'���I;��Oy�JS6 Z�vM� ���&�?T��a�a�;5(���u�;�IR�}18�=����YG�.�{�s���� ��j�PJ�f���xZ�n�V��? ��`Q�ޖ�\/`�b䂳ܼ�ٍ(�?P2P�<��'�]q�y�pGB
��S��y���ko�����=zB�d�w���c�wg���|ު����A;p'��|̘�sw��~�B;�Qp�V�?���u=M���Β�li�GO��ץ�dV�xѪ�u��F���n_U����E'�B��́��6L����U�MR^nT�D�k�1F2���e(Y����̟�A�7RcS�L�1v_v��o��:+/;=��q�	�h#�#I����L�K���X��l]���d�!oն�miP��8Qn"\['��k
8�a5+���xn��PH���6��[�kL8+��4���R�F�$�*�G�e�b��DZM7����N_	�k��&Pr�Y��0/#�o���h
M9]��b���?G3��V,62���T����T�p��nB3~9��e��~k!�v�n�^N&���r�r\ 9�4smq�ytf���$��|靀�=�&#Ev��~�,Z!��DOA���KDB��<��6��7|m����m���A#Ze�|�N2l*xh�9�a��1������h��կbZ�yA�*�j��3HW��"�L�]e�C�ٰ��ذhI��������� �#,p�Ԓ�	�>tV� ���(9{�-�6P?$��j��So�sI-~9ib,MUR��AS����{I	OJ.�J�<1AA�dd|�Dj׫��&�H|����_���[{>cB�;���aH��,��}v��~^�;#ַ_]Q���GT��4kK!9F4!i�C��,#I���h�tܾ���{"�0��m��㳡r�m_��i���$��M�����C�5���{��"�NW!;��A%GQT��{�\�뤳�J�n����F� E\��2|�I���_�������e>�o�ܮ^��=]���ˤ�T�y����^ꍚ�"y�U]��h	W"6X�d�'��>Â`���w��J
+R�<8�M�c�|��>U<�R��p���%�f.FY�տ^_`���x��I��"�7r�8��1�_d-	�QEAg�l`;l��b���\~��/e���+��ɢ@�d���m|O ��9��Ԋڍj����B����s���OE
����������=4�r�J�(r�N�-=)m_˫0=�i�E�'�0r��0[@����o���b�I&����k�CJ�0.�_����h��7�VG싰\S���?��e+�D����V{��W�ڄ�XENVb<�JF���~��'y�q'I�w�o�m���E�<����,��,�c��f!�yE�:w�b��J3�������m��?>����)�h�-���f�4��D���I\��χ�s��:y���O���4�4�	�N0	���pE��3���2�x�b�#�P���O'0r#J�"ӕbξX�S/ �{����+�Y��%���T-:
$�	�ؖ�r��M+�-��os$�o���m��fw[�$A^��I�5����p����y9��Z�v�2݄G���\҄���t+�R31����"�pU��ɬ�F����ﲽ���G�|���0�l��UU�	�M����3�uBPq(�g�]|� r�[7��l�?2����aoThRB�Ssr��=����?�
'��K�Vqz�nzܿ�C~�6���vmؤ�϶�)΢�:C�8�ũ��٠p�tCc�O����g�~ׂ�WGR(���9{Bc5.�p��\2
~Ph�ab��@�S�ҏ%�nE"��/� ׁ��1�X�ʙ0?�N���>�!i�iE�� �P�����[���)��"{4�sU;Y�'6R7 `�d���&�m��6�Y��m�GI��g����������>9;��[�3�)[��\�k������W��T��V�Gg���qv�gB��2C��
�ݙ�'����ĥ'�H�&6��~"����*�sf�@�����Ttq�ow6Xr�� ��S��c�>��TW. �C�@�!�d�;��r9T�L�q�ꁔ���Y��g(l�P��������>�kEm\~E��$i43�e���H��f0kIIťY��C���G=�0� ����˜�+E��W��?���4�B7�>�F&Ug)o�����QM�(P��W�i��N/_�@0m?9��|�*k���XҀ��͑��hf��t0i��M�v��a�J(�%5�+��VP�m�"-�YUo��Jp�G}S���.���$m�"'�aj�UP4���3�~��������mZ "�'�l�uBV���ο7p�C]>�CI{����������[D�dgD�Z�a)d��Q���fs�]v~w>�&�H7p��vE�VJ�L��hl/�E�r�	�����e���i ��T�;�y���+� �>��Ƃ�;������tB�	�@4� ��Y6M���v��؜5m_k�+b�v#���ߔ3��ק������1+J�@�d௞ ��\~����_oçkPr#�cC-�v ���:T	���`���q5��7�����ˮa���,�/,S�q���2`������������,�A�k� G��C�Ԅ�B� ^��vZ��*���M0RR���E[��|Pheq"s�Г����u�����R]ה�]ں������{E��_7��o�Eܜz�����❖�钅{�R�v�ȯ2�|f]>j��F<�o� !u`%tX%ҷ�s�@��HY�ǿ$���Њ������|��\�󾯥r��������l*.���ȅ�<zo���먪�$�W/it�(�*�o�7�ʻAvڇ���쮛�k]��0|�S�\���.�4��+d1$. f�\2$V=��e�`Z5���n���ٻ�a�O���
�L��l� �@U"�Q�Ct����|�yɕd�ѱ�:X�@�o�����_�k�%��Y��& P���=��Wnl�4�]	���IF���vh��B�GY	C&蝈֪�:�o�5�]Q릺2\��-@��(+L�U�}P7�N�7�������s��J�9{7������t$���Twr�-2�4�aj8CIX����c������������!�����
\���9%b��mkp�.fO+2s��ۖb`�C
Y��������_��N��}c���R��]��Ǡ6�0��$|_��׉���{�7�%��rO:g��;TCx�E޿w�,��\T�:Y\r�R�e�J��-������l��I�t��}��,�_��c��TY}�+c�.~����ƕo�rv%x>��K�W+ȀCм*������+�~�P���@Mu�ZWͅZ�:2�oQ�;�m�-#�˶��k��r#\��~QXIut�8�{�����b*��NɍUw!�T���(zτ���"
q��x4���Ufԝ�:r3�9̛��&	�m쭡�h�V@����˝�,��_x+\�ՠ�Ϛ+t��Yg=z���&�"�t_�|_�SS73��<�ȵy������	-����L4�M�����Å��,>*�������~\��ӽ�`�&�G^�1�����s��Q(>�%i�G�l����jh��k:�j��10�Hex��㾐�0���gPb��ڹ0��;)�mc�~+ڜ4���'��:.�j���,r��;ӥ;Ȧ�[�٭�F����h�a
9��W���Q�=�:��K����-�Q�$6�c	���D7��r���m�K���D0kf]{��)�i���;��b����W�\<|̎ނ��Ml�,���>
+*@�U�2�5��k2;���;5�����j���f!�0>m�8����U@P.Vz�63�d�]�q58b�s�ac��Ԗaԡ2r�ӧ+{{�MT��<.0u0�އ�3��Xq�\A���2]���x]0��%��)�\G]��ӣ��A�}���9���q�uwW�rb
2K��-E�N�Z�No/�t�}_#�(��b�ej��:�����#����u����f`��l���xM���%�`�z�v]�O᣺l�f�
8�TJ4�����,8��o��Ek����T�K^�H����kh�X;��[ů�n��b`3n:g%���%���X�A�'?��a�xB�� �X��ѧra~n%8���]�gBA����,�y�$Sa�.�4Q���1�!�[^�#��k��_��xp�%���]Dl	72�_6��,
2') =�$�v�6(uK��IR�C�@���/���\6#��U��I�S���\�"G���d��s�i�Z=��ui&�� 8�3�N�y�Tvj�k�&�!� O�� �i"�tY����~��
�Q�s :���G,=�J+ְԛ9��6QD+�
J+쑟&�$@��p�Q�s1���}��#��m/��fEpruG��a#���t(��,W�Q��Ϧ@�]o!���$t�P�K
�!��U<���V��TŽtk	-��z-�/b���<>!�:
ر,�%g�}Aq-��	/�q�9�7P��p�y�тY�S��	�������N�f��~��oQ����h��ô��Jrx<K��Y�@POC��	9^�t	[�6��x�f��*��#Iz}�@�>�k�ʀXB�J]�]�&��$��Yy9ti�dh9S���7s� w[�<��&#���	�n~�#���\��%VJ����&�x�ŏvR���r�+M]�{`Ӄ�a��'8�uKx�}B�rX#�IK���zZ��8�X���(I�c��z]K�ގN.��m���iOlV�5���_ O�.����o��g�Jx��V��iMCi�x�B�tM���)XS��k���`&o#` 2����ܵ���_���s�ߴ��je}�)d���a�9�|C�&��0 �?}�|��֌*���Yγu��;���Goa��#�Bw���|��/�(������~�-?���5���-M�K� N=��	 ���?��ܽ(>�Y�؎��E%*Y�<A�� ߋ����ݘv�^�U��$��+����9�A�+R��DE�^�"�Ò(n�::H�%�' �%�r�*�!�ن�*�#�	ʫ	��UZH��.1EN�����`�@�ਵ /�;r�4Q�%Ӫ$4t�}�S�m/���.�u���K�J�#h�c���X�]G����N�=��ڊ�]A=�_��mf3R;��ȗŠ�[��&�r%�1^B�"�jNnEy�ϣ�<�r/���cM���C4�"�.A�3$��{������l?���_!N,�"0zg�yn��ŭ읟�x��3p:-r����q�Y��A���y��j)$"���<8;���v�5���	hBh��O�o ����e�ؤX�^q��N���	���v ���u�3�����+K��[�7%��Xn�DB6G�y��l@fV2z�m���v��`����\B7K,�tM?R>bF�qw'�&
��+$�N |��O^u��5=������`�����H���J6���Y%N(�z�Y���L��iPP}�p,P��_w#&<U�����[��U5X.� ��2�i����0�c��:��
�P�li.�����E^�ߏ#��MrW-YJ�d�;�q�_W��N"2��iMG<��J�
��o���T9�Չ�X�J������ {l����WTfI�!r�2���?%=s��Q�!�l��sl�h��y+o�v�Š�6=[�<���=ݔ=�`�����,�����y�_�3w
������N�u�ɢe�Ӱ��N}����_t�2�EoI^���O��aW�(�ñj�9ax�����{�z��=kh=�����6�&���j|��]�o��SF�`B��3��F�\���U�T�o�+��ֽr�Z����V8���Y��tW&�|�1§����%K[TȦ�.c��7�&l�cT.PIWU�~����3�m<�(/���h�����3�L<�xo�:*��K� �����=pϑ�۵�gu���@�Ό�ҥ�ق'�=�.o�ÕM��B�
�5�F ��i����Nw��,&i�X�B�qtL��X�?\qu݆���:�p��ٸԽ��zu
r:(f������%P�u��9;�J�R8��
:����E�|?rc�P����$e�v6�oQс�}Y�K)���Yq��xП\�˄�u����fߨN�g}��{[f�Z_ϐ�{�� gN�&�;tr�������Gi]�\K�5ܸ�6��u7�r�(��E�&��Å.��i���f8��BOm���B�0);خ�F+9�̀�����Y�J8O#��Х��%|��0�2*?d%�&)���^Tyc	q�����$���;bk*�?�J�����[��Ƥb	^Y���Kݏ�j���	�'F@'������ω��LO��o�G{�2f��q��9h�暀���d|m�W!H�+�5y�j����?�B�#XZ0ؤzx�I���^%�?T�"޹�0��%�v�E��
n$��]���t%�VE�2b^/
x�uvM 		|�	;��+������G���U�?��v^T�0M�;�$�K��9g���Zv83d�� �g\D�	4B%�Ek�a�t�~�A�P��r�<��kX~}�W�� Cs˪�Y��� #�]��ʖr�g�밒���ڏ�+!��F�����W�E*U0�������Cj��m�}0�;��������d��f��_��܊i��v��_AA�F-7B'lm�s���׶�:�(}�HЙ�w�q�LaF!1K#�y<Xl���i�@sv��\�лi&���E��%;b>��MS`ad��U���Yhß�N	��'�d�	��9	�Z�<RDN�{�7a	��/(�6�u��ci�>e@Y?�{�@��cׅ�� wr+�T��A+0�a\8~kd�=��D���ܫ�ٻ���(�pJ9�g���ag]Ô�³��Y��VE���l$���G�f�gW��v�`]/8]��� :�����1����E����lt>�ʃC����#��u"o�<��~�G�Y"ݟ�����[���5��/��>HZ�n�����t7���
�&��m��QVZR���,�L
��;�G���!�n�ٶ��8�KFU�Ԙ�Dx(�P��~V8�9@r�9>;�c�u�f��"�@ang���]�w�㙟��cf��mf^W?�Fbe��"I��NO�GKW�/L��A���G��{��`����f�	�@�*�ٙF']��>��Z)(���}p'ez��R���`�����ػxH��%��*F���c����4w���^��#����K-l�1=����"Zk�v����E�	e�������!̒=��e���5ǜY�cNr�K�uy��/]�7�uV��y�H��=�l�#��N�h��''}e�DO�9���:>���WH:���ʅ�~�֜Lz؆�NK��}oc��V����~���z��?C��1К��",Է�L�Ut�]V�\c�=3�f+ľ��C��Cb$��!�~���T�Mp�|�â,I[?���wD��� dZf���0���*�����pɍ�{6�6L�X�4�z���N���r'���RS�8�w�~�i�L�nOT�w��cn��"鏝0�� �\&xs�P��⢱/l����>Q��y|G��k��~ogӌ�������ja�%c��&Ɋ.���0�K�h�)a����GS��S{̀�߹#�_����#in1;t���)���g��M�S�lt�Du�">G�MѢL�?"l������#G޵�$
����X|YZ�x�JH��p�8Z��&ؠT+�_$uۦ���"� �tQ�&6q�و$G�"��a��YT�ч.��q�9�X������qh{҂o���-��%-oB4������� C�ޥ���	�4�����X%��C�K!�D;��7�)e_d��Q�Hp���1q*��Ȁ�ϊ�{(�I��}�0���O�V��� "�_���n7�V��rR�i�7�#R9k���6���|Q�����>�j{��D7Z�5��J�a��p{��M"F2�_�Wl��!��cT[K�$(-{قy��^wps�$�4�T�M9i�9.3?!�g��3�3-���gV���(��|~d�F8�1`o�/i%l1�8-�ֶ�*?�a��Ab}݅��`��ZRhj��L�*��m@y�~t:{�c������;G0������C�GGjV-����h�+s����_���y{WH��?林���'�W�;���J	Ē�BY\�v���F܁����Ge�w�Y�!Ln��C:w�<�S�)����_}]�*�\ѯÐ��dr�9�a���FS�4pe��f��{��Xq$�n���^�mЯO���*t�Ю[0Xb��Qu�JGˀ8�^�$�[�[ū��;Ph먊��
�~!�|����U�(`S�)�����oy�HO�}����YFj�*_�y��z8�_e�]&���a���W��n�1jz[�t�,L�R�1iq�����]:�� �G>Q�S�`�M��V�|��5e�
=U���Udf�����)�F��Ƥۏ�=��R"����L�.�_I�rt��/+
�h9�t �c�6�Q�R�`������GBtS���KAsq�cf�cP�{0����b�\�P�d4Syj� Z�L��r��/��9��� O�w��j1�b�[w�V\�3�Z�n�ԣP�wZ�}tm�g��^f�;ZN��G�gN#���EL��a1�m�����~ ���~�g���.XՋn0��^����5`���7��V�%�f1W��Wv��齵�c��n�h�8|� a��fSA}�M|P"��r���A��$��+�(��r ������GԢt�;�%����01�����F2(��9N���?_��Mg�9��@��A~�V�o�śz:������)��G��~��8W{�x���,����9=%�R�_CM�|��݅b7���fȠw&�xu�8���SCߏ��_K:c�\=�g�l��2h*؊Z�\�����C�"�V���p�e_�r�0^zo%���2��3^��ߩ4a;ʳ�P��2}�Cj!Q���ȸH�j�^��0�n��/��K�'��w�u�"}*=�$�8�X��M烶� ]6ª�I4�ur���MpS���scџ���%y���^�\�^5h�-?aX�����E��qȡ�s���J��Tɧ[x��x%�C~7wu�X�B �'�#f3�f(��y��{�����ūQ3�;Z�?�;�����qu�4e����`�5�;��}�S��!�tn�Jxm�Ó��!}��hy��BƋTm��{�ň��R�y�2P�ݤQ&:gt�O���VX�H�0q�.�ד�p�1����Gc�y_fec�\��i��gw�������S��R��/�>|c
=>����	�}�E��>-�����dl�0րG��?9��7
 �����q��b�,�I��5s*̦�1����ga��ь�J�v���l�2�2�;�A��$l��j^kR�]s��{�F�-cc@���Q�D�tt�-��p/A�I
W�<�}���hu��H��E�3��8�寰��p)�[g��A1�p��. ��b�q��ݢ�\��ێ��Z���M�ǥ:�	I>/�&���fc�g,�快����ؼ�҄*�)� �h6��l��u�|����'���+a�#�;;��s�-V��%/�+տgL�mƮ������0��&�&A�K`^^� �?�A�x�4�}8Q�\Wb��:�ٔ�#:��oO���á5�&,\�Ku7�PFa������|B)^y� \���n�%�e�~I�T���Օ���M�B=jh+C�BA��Ō�m{,/Kߵ�yҎ+��QƏ�>��]O���&�m�Lc�w3��$A��̺�gt�<��B�"_���8����:��f�$��XQq}����h� <���S�#q�A<g�
c����?���w��I�w8\u�����]:λ=����>�IC�^�6�ȶ��n�>�.�5h~W�E]�I�y(�m���k'l��N%����hFN �d�TEh{aXv���]3�TE�*MF�����gr\�������G^W��&�x�E��亜I��V�	����ӂ�{P�����c�N�c��&��A8;�o)��7[2f@��w$�*�!��I��f�k�w��׭�l	��8x ��]���`���y�sʠ�)��cEr�:�8vRi��	�S)�ˑ@����|��>�N�l����{��&Ϩ+����-D���Z�暚���͎��=_��o����@eţ��tY�&��J������*.�j2l�Ӗ���@��~$��hZ�c�Rf=�m��������WӢ�.i�}�|�6o�OW����H����8)5W[�L,f�"-x�c ��#Zl��g�D�����'{��:4�l�X�c�	�)�Zô��Lؔ�S�9ͿPj�!��-�__��Ǻ:�`���:�Z^�@I�m3ǥ8����\P��YZ[ϫS�m��Ң�u=� �[���%3�쑄Jd� ����d9\��4��ٜ���}��ݥ�40�^2��lr��}lHN[|adj.�Ǆ�r�h٣��l����خ�.>��sQ �c/�PMh���c6�Qѵ4Z>ϰv�2��%�y/�Fw=D�"g`�`R��W�Ӫ�ށ?z�Ni5�Z�=�Ŵ�4�4 �|ᔄu� �M����q4�-ut��Z;�ZiB��dQ!�X��Tl���q�uAz�.5e9AWbeC>���u�/߲��h�#fͼ6�� z�-���~B���I��?��l��h�V#�=��y�D���񯳴���0��[����-�6��v��dZ�h�����ؐ��#�=�|�b/��F/���~��� ��}��u]���X��~���_x�'��2t'.�����"7N��m��[/�5(Lƛ�M�:�F)�<��x�IE��~�lP�!ߟ��h"g�:��p�.��F���tGu<2�%Z��{�#B�̄Ei`��q|����o$�����@<� 'Q޲Gf��z-����WvC����	�D�v��ٱ�U�\��T��HˢR-��~;�(>�I7�p.���z�D`�9,H�y��"%�K�R�wK���xM��|8�~�S|:z�;������3m��xs1�#΃�[X��F���殍�IrPRm�ᙳf?
�$%|�"��Ƕ��3�C��J���`I@[��
>�U�q���溤E}O��}v�t�#B���s�N�:�K�T��o�H����.�ӌ�'(N,�eC䵔`z.0���Z�/��������7���j��)�����h��yq�[e!����sT�P�SAu͗�>�n�N�)�'S�R��m��K�*��p�����$�;�H#�J�G�������
���dA�����˿ܙ�|��ֲug���h�6�U��=�gW���m��J�>K�j�����{FF4�Q�8Y�|���#5��m'�t���
�it}�X,�'
��_3�Zw�蔘����f�n�H�oh�o�C�[�;c �Z�>��*;8�hFw��S'�Dm�-Ct)�c6����@)TH�-�X�q�{�}��=t2%Y(_�r͖
V���iY���g�ݥ ��3t�����i�B�2 02Z�[שESh��6��n���8J��0�CB�β��%��@����I��ELwf;zִ�(4�/R!s���$y�W�K��ܬ�x3�#	��7G�_�PN]r�Q��=�~��Z��L���̼�B���vv�����>m�#,kOm���<1��=�$���m�,��Y������ץFע���#K?q��|�H �WI����h�`�d���� ������L.�6�g'��S2L�(l���Yx�;�z3v`����h7t�h��[��V�{����
Q�Τ���.||#w{�pPˬ�F�꼩7P.Fd�<���uҍ��;�`��s�0p�l���L��1k�.*A>�x�С�`u�
�(�:b�fe�Q�&� h�������a���}�7E(N?;7Soe&�'��������}�d뉒���bm��2�AsL��5��}���p���:�z��?�h9�+�*fṾ�T$a�f9z(8Y�D����Q��B�����_;+x�o��\2�2��/(����EC�ML���P�`������3�����"��iY��yej���]��]SQ���	��I�pKlC��ć��f����t�*����@��ZR����!X�:��pΐme�^���C��욃��:���L��\%,"�Y���sb�Љop*FC{U��H�l�җ%�zr�hF MłPfz�P��{�R�E���!l���e<�oj��LP%<O�\!Ȅ��r�؀�F���_�V��Aǳ�V>�{��H3��8I?c���JSy����T�x�Ҹ�Ԉ�Y}��E�������?h�d���~��E�\n��s(�aP�3+eE���O��lyr����0|����<�E�R��K�ŭj�7��I�)��Ua��8<GY5d+e�sܱ,͠�4�T�>�JԐ������'@�%�,Nv�9�fEvZ7�(
��kP��q�l�����<4�.[���s�����`������rjRr�/Ӹ��͸֠�� ]���Am]=^:�,�ޙ~	[*nK675�`]����������jPw��ҡS���̨.|�z�������C�BIR���{�h�I+�Ϩl�Z���R�����ܜJt=�;�h`���P7��Y�vK#BG2=*Xˇ���{�=J���oU�y�>����Y@�����u��l��^��-���D�r�n�	�E��-���{���P�V�����ugmb���d{FN�^%]J%A�{�7 !����NI����B�=M��^�)��qlK1m���s�VQ�9!�H�siA_�`j�1�F�t�4�s�r�V��ؘ?��xֿ��|G�9��s&�o��軪�L/1�J(#h��^)Ǉ�f(F�%�Z��l.�Zz�;fzW�ݕ����CK������58D��G^wE1d�`�W�՛�����I�V`��3�輶;�t��h*_!�����%`~ 
�PVuH?BQsy.��V`&�qx,H�FQm���@���X��;�s��7�v�o@$r%BEC��!�b��$�
��c�F �ݙ��L,R�/��A�+O��m����-f��(�ex6nn�&����_:�cw��G��N2���3�����|Ķ�g0��Lx)m���T�)@�� ��l����k`b����Sݜ1%&�IJסۅ���Z��;��ٚ�[��kZ�/+%�v����~�S���#�WpYjL�ej�F-bo���u�kgh�P)XT�,/��{DJ��t���}���ϊ_9��h4���ZqT�ޟ�X�[�뱄}�̉���S@��o���x�&1�����O�m/�>I��Ŷ�[�(����jW��3�F��򆗑4D�ޫՈ�,ۺ�\����rYdS�?�Cb��22h3�Q�J����i�6�2ᑮ���d4�cW5�m����A8&��˝�� ��l�����i�/g:6gF_�<�[�[F�1���Yw���d��Q����ꖊ���%��:Q!68=v��2=��E�o�M�>	�0�7�#v��<{�8P~�|	�##.{F�3d�(g5|���?ܤ0�F��K���C�:�v���p|ME��<�$5��ĒE��7���ǆc�c�]�:.�u���z� k������Y긶S��t�rH.�D�ﴧ�G�F��-p�&�	�y4���Re�bp菜�����Y��Z����등��cW�X�Ģ��{/vPM��W�RqG�2���c9�|��!��N0ܪI��`ݘM�Q�rl#� y�:4+5��r�
i�ϥ �8�]�%����K�)"+Ys,����"��ه�.]�9>�<1���Aj�bHv�1����M��QJ�W��l�4�a���{j��R�5k���z�o������-c�iI3vOόşx���C�{�$93�U ��m���]ͱ����qJ�����|�H�~��T��Nĝ����f�*�]��!ϙ=�J�q%C���I|�K�'Ë�:�B�k�y�l�?jn�I`���F)� �!���%�Vb6k�b��9��x_���{�ٽN뺭��LJ m���Xa�g�/��[Y-�$�g5Yd��B�|
� oo��s�\�en���럵�+��D1��M�Sȓ
�5c�%�*.�罜�C1�-OfQߛ�:c:�L?��=�>�����,����^���!W��|f��Bg~�<M�~猝���Mu=%ʒ.�����]�$)c�鮼�h����Qw�X[��髛2��m�A8k�j�'#m=?� V"���8�S��K�r�[SJ���١�2�JF�*�{�V�
a;ߏ��
Lu3j�	&Z`-����祄.����W��iؘ*zA.�����E�\.c$�����q=�>��=��V1W�6}��k�^���*�'�V�S��,;=$�~9��A��$�5�NY��J��V26��6c�D|�㶇��2�D�dpA�Q�Vs�I�ƛ�-������|�.X��-<��*�j^ ��]t�&%��֡"��D�-F}�c=ĳ�ٴ��c���B�>7B�sY��@��J�9Y�y�T ��8Ŧ��8��R�9t˚���+k10�&��xF��?Q.�����t����@��(NIf����W�h�xDw>ּ�~E�3�l�]��k��1w�`o	p̡���/}H�w�{�ig�`;�(����7jO��;/-�\�`�K�l^�� e����W����N�r�y�W��?���5�4��g}|�ڍ鄜���h?M[r5c���8{kp�\^%R>�Qfy
��Xj�Q����-���b׫�E�!��O�׿i�q���rT��H����f��ѥC�4��7J3\'2��k�a���}����9G�Q�ߙ�ɠuL�&��?�+�L[�9�_�����
q����FQ]|,!~�46~}�x�5�I,�}���rD<_���.�R�Ī{unh����P��PP{�@ �Z��+�����2�#���L���Bt	r�RI�${�z�蘐�����U&��1ѯ�s3
�*�q���� ���@և�!+VTWQ,Ӫ�13�r����~ȄʸK{۰{k�����T<�p<�,#�=b2k�ޠD�U�Ý�6�_�I�PP*@����Ӝw��*��c��-=�a,�C j�-?פ_��/�^]D+R,��ޫ�����n�*��V��Z�$0����\�E��g�'�-B�qZ�wN�ee_!9a��a��Ȳ����^Kd�z��d@:��+�������L¼�{���I �ﾃ�畛�r?�.�!����3q���[-wD5�|SW�7o��U��R~� D�F�a'�p]Œ#*����/��uSn}͚����3�1:��κ�Y����L>>�8�^�a
t����P!�^� �������n�}�-s�ptĳ���Mz�O"�����a�0�F��	��z��h;�Gi>��@VS�����E�(WT�n=��g�޷^�9��4���1�s.qƎ��6����l��~�s.��E�>I�0�6�pט�q�����0?c�0/�p�B�C+�Ww0~�6�W�~��W�N`�-Fל�ƋV��c#�Mg�����9M��s����y
ۜȀ�Ŗ+�}0Xmr���i�z3����|��ɰ)��7^�{��a��t�gk�����:c��i�;Sg����E�"��c4�+�(�*��ѭ��r���;�r&~S��&����i6��F���s��բ	��C��rE��ŉ��N�Dm�0����| BQ���F$���$�M3� ��_%Zt��u����s�B0����
f��Q\�tD�,�U�j�O�N�%F.Ck?ۮ�h����9�"Z$D\��j���{�hn��(�j	�Xܥ{�%P~j&f���zHށ��K��`·�X�P���cC��H�ߡ��r�{6rtY}1���S��7�&��i47�J�uw�5WT��]t(y*��
M�m�{2#_�F��P���_���h[~j�@�)�L<��ʯ���=~��vރ��q"x1A%�. �5��h��c"���D�*6�� �M��y�FZ��h?�p/	����i���Y/I�:��[��O����R/�,R�\�#5�)�A�ջ�քO%?u&�ק����?`��I�#��'T��X�+x����¶�4��X!c��
tn#|X{��� ��'�@߮u��U
~ch�ꩄ��1d�%�� �!��_�:c��Ϸ�ނ�w���,1,�cBhS7C��:�1/�r��zx����/TV:�,��9p�#�T1�{��)��N��CM�T.�+�'Ō:�����{ฮ�����+V6���3Ǭ�JX��?�_�I6�����/�l�C����9[㬕
1�ָG��.�Lj����h�A��}-��diaS�Q��%m��K' ������y~���k�u���͒��X�u>l����s��[ړN��tB��l\v�+�5��m��0�b�5���N�?�N2��Тf��ܪ��@ ��1"��Km0H��{���ks�)t��G��:̣�T�6I�W�4o�TO]�� y�S�tP�B (��_6L�N��,�!ߛr�A��ŋ|�4��W00J�����Q�S�+>-�AR/z ���M���7��`�N�m�b�όNe��w	��ݾe�CGL�8�m��i�QΟhS�slqg$3-�˰���)i����U��1�3�yY�V�K�/\��=�1@���>�7A�pd�^�z�C�	v?�	�^ 5�$�0o���9�ّ�ލ����\ҳ�������՚v8h�3&o���_Ӽ=�?zl���KFϨI����6�{�G�	 �-���҆�
U<x�C���bZ�P�3E�K�2|����8Vp%3RhD�Μ�L
����Z�ߔK�KT̙�k(������\3�F�K�ר�=����r��n9i�""�Y����8���E��0*���-:�gTO�.B�"!{���9�f � �1�w\�='�b����I�������W#��Uu�0�$���s�+�֞7�Ϧ�F|�)� 9���kNL��uq�j�C��b25߸h?�a��עw�t�H��2��@{+�Ļ��+\�`Gփ�<r�����M�RA��u,Q�_���r�[]�V�]�L��3Cg�X v�U����s�J	�T}�ւ�3L��Ә*�A�׻�W���p"^�"l@�|y�Ѣ�E<���,�~J"�������%# �B��-����\�����B�T�${Z��U@�w���8��XS6s�!�(�Q4(�嗧_5sO�V�ԜA틯�K��oJ�o�R��T���j���O�!��s�Zy�s|5��?���)6��"�T�Z�_Mf�D���C�V��qЫӵ����`]�_�B4c��G	7yh�����p3^g	�%��}<{��ca���vtێ?'u���Z��y�V��n5#��+�{�Wm����u�UH`b�fG�J7F��dsi��%{�õ�����݆�
x^`r	J{>qc��&
�������r���E��5�ZaP"�������.R�/bqv»���.��D��Jhk��A�\��\
���u���6�O�L��H�����M~���a����<���<�j�n=�z�zgKd	!,��5ttB��}gw�{_�3�cB��<�M�dG���'�L=x���T�����E+�Mu�>����T.ׄ�(���!�s����qzB��V�n&�=/檐��l-~`U��f���!�`S�ٷ���LF��5��B�f��:)��(���)��@��2�V?/-0������C�q������/"��M�w4�D��cXe��iU��^�vu��ZH��m�^��O��޾����|��ѱ��G*F��>>DͶ�6S�U�F�L<�!@젨��%��bzҪG9��b�I�_,�S����������s�	����2��UT��2l�������0���`��d��P>�����c:yh�w�L|wA�@��!�A�[V ��������Z4ۂ��� _]27�J���O��^��6�b(���7�[�h��t]j�	i4t
K/�5�nRF�c�T�j���Y���mc��%U)���"ׯ���̜#��(��$fi� ?Sj����`3�j"�H����PU�.}��T'�"�L�z��������7��Jkd[��iX ؼD�q��X�y�U<j�tZ�P$�P(�Y�q�\�?%�B�T"�l���I&/���>���U�ԍ�]�!�TƯ��gWI<��>3���+�:u�_��g�, �<�Bѿ�����z�9+��@ML#En�|�][���X��4?�m�Յ�;��U��s�M�@ɨ�=o��@��0��8���3�ĵ�p�I���)������U������u58����PGI��ƨkM�����׮��D���c�uڪ&�0S�\��xSf�� nBv���ڻ�KF��M��"	6�:���?|�c��$�"��n�a?�d^�f�/�G��:�۵��3<��z.cI�c�>�h�Z�%�=� �+C�"b_�z�~C�zuS� ���d��-R| ��"�����L���`���+*�
3	��D`�HSB&�.Ù�Ν)��(�;��9&�L|�^�v�Kb�1�M������H�-9��CċX#���7|n��o���)N���PAXE�@��B�l���(�ڝ�-X�(�_��C~�.w�7zQ�ﲓ��c1��L��b��f��rZˍ�aAu+���a���ݮ��u�3�Ql��0�*���`qˑ��:h[m1Yd
�L'p���,��L����Q��W���2�6D�Z~R ���\�.��͆^O�L�Y�������o���*e4f�1��Gxr��eږ[�m��bq�L��;eq*N�r��ZV6"W�>z��W�s(�W!�bh5݌�_��ڊw���/��z�>d2 '�H���!�I�z�Y(�!XB}�&�{[B�b��у"|C���H�d�\fYU���BNW6C�+M��|�qS^w�<�"��E�[o�}g7CI�֚;Y�b:_{i<��z�]S�͌8&�.!���h��"�����ĵ��*�W�^��З�ҌW!���C�Vt_Sd��:�&m;�q6�.��)�v%�<%�˄��mGc�v�����tA]Qq���FfQC�\*\�A��f�d��`òo��&/���X.{��Xᷥ3�ľ��d����/�h$$r�?�����Ũ;^3E�t�S!{ύ ��=2��,��R�R�mZ�L(�C�F�a�y��������FŲ�zʭn���8��(���C/e�];�������S6C��%�"u�b́|���&#z��RJ�<Hl@6��d���ҟ�Rkl��0Y���?;�XW(��e��EB'o��a�U�O����"��	5���{|Hɼ��t��Ѧ���x�V�B�����Y�@qW���P� �>6��J�*��
F�W�&.(��l�f�wPÑ�����o�2�٨��p��=��΄89q����y,� ܮy���R����=����o�0��U}�)�"��k|`���/(�Б��Ɯ���A����un}�
�o���6�=OU����4�Q ���r؆ޭ�в
H$A���N0ڋ5�-{��Voc�T�M�(̔^�Q�n�]����V���	��s@v5Ǉ��csv����)g�fր9������+��/Ԭ�
߷�Dr�@�u8�8b�+/[u����r�I[ݒo�,�BZz0DH
��Z�����Q��u�M��o=�z,u�%��g{lq�55��p�;����f�[*/�H�M��H�ˡg(�I�w���X;S�b�-��1���+JerY�}E?�� j���r�"��N�:ڹK��;�P��U�1��ˋǈ_Ӆ�X�R��@�1�Nh����.Z�s�_6�݈��'��\8.35����Q�m��@ҁ%PtCk1��l�ؕ�`�kY>u ���5�]��&���Y��?�rx�o~L�S���Y1R��ӵ�S�Q�J���I�o��h�h�A�g�l\Dө�~�BAɋ�ν��� q4?EL:a�#Zפ��PΞ��.Y�\���D��~���� ܤCh�#�Qɣ��G�VG�={i��/%\���}s���FX��2V+)��!���d�\HX���!��:��5�~3�u9&�Qէ�N��G�R/�^��)�r�O��s���o?'|�b�Q5��.��?V��� �`�%�LM�mC+,�$�lcz�$s�}����z�{ƺ����ꤟ����_
�C�{�٫d����s��/.3u�(J���& ��gtA�u-��\�4�n���1"&�?Gﳭ`�N�*befZ��u3��O}W5�U0ОՐ��_����fPVՋs�G��k���[���F���n��<v%�ՏBAQ.|؏��hɅY�=㡜��U�v*ӓ1=���"ka0
 �\���Gњ�k�W�0%7U�Q��Ш���]���#b}D/���=�n�b=��V��\F/r�s��٥$T��n�0ܒy�����`ڻ>/�Z�Cy���@)؍�8{p��*�C��'r��YZ�
�Q�b�j��`3��g"O�+������*{4X�Me�(��q�LQH�\_ERH��}:D6�8I�8��(ƫ��iށ �d�	S0E�̥-~so��l��G�bB�N5���j�Ř��;��r�\�����p[0 ��)pQ膻�b3�E)�<dMԦ�/�ҝ�X�_g`H}���ǬK/�b��<�Nq"�VP���ao�tP�]K����Bt���6ΑG��X�˻39bRv��������XKgf�[H�T��N��& b>�A�~+.��ↁГ^Y���g�nÄ�W�l1�4�GR�6�d�0�%z�3.��f���wg ;��I��i�nzH��{o��p�,���������x#%΋���p��jYሉ>T/��|��{���ވr8��ھ��r�#�|��Ň�(Bk��ׂ� �(�z��{���[��=r�{�V"a��ZH��9���(��-�.�{}Q#V��'����[�"�i�5t��C��?�P�ޘ���6�K�
���$wSw�J���h�잏at��º}��F�U�����jz�R� d~���\�Y6ߎdY�@yKy���4�[�Xc�/<�q���3B,B	�1���[gm�+�a�Bb׋�g7N���∋��h���CW?����E"H��+�p���٣�������n�U:�ln0U�,@���0�|��L�_��-�q����Q���fy*p��D�H�t�f+Ѽ�9m�/>����4ٻ�$�ƚ�>)MH˛�9G-ʙ�[i����9vң�QW-���#�Ś���a>R�o��e
��)��~��X 4@l����8 �e��\��7{7�0�{q�7a�ĝ�&���6;�5��Ұ�ٻ(7�>&b#d@0�@}�	�4��w'"e��9��d(����)�
m��[P��^��h�ƈ�����l�!v�)�{����6&�h��%A�D���s�VbgB>(�-(�t��H��;)2�������.��G�OW��R��oXb0�^J��-*���R*`9ui���Ć���r��T�v��/"�i���v����ږ ��?W������bPs��v͍��`��ʶ�*�!�{��/�Wc���JPMa�������:����ܭd4����25�(\u�P��Z.Ծ��%�l>b��⒚�e�Q~��D���`�)(�.t�7W(�%u��'`�Ӻ)�rRV �H�mv�9FmvM#��_J]��'�A��,=���ݝ���ʪo���u��HJC�6������7n�Â9ԩ��ݷ#!�i��<0�,]h0��e�\��Rϯ�{T9I�iz�ޘH�BM�O%�:��0�%kۑ|S�0J���!�c^=�Rq|�P�K2�荂�g�L-�D�*�Sx��n��e&)�.�u�a�W@��ļ���騿Ls�2�]���0�����u걉ge!�ކ �EԼig��$�����-&�r����N��G�o�Pj�О�.X#[·V��Qg����e��%�@(��o��Թ���8=2���xui�����G��wY�n 0:�k��	���ۍ5?Z�}�ѽ1�ʦ�]L�R�hĹ9Ǜ��}.�t���r;zK��h|����D�Dp��y��8*7�e缁��CU�gw�kV���6�\Au,*t���{J�1�*?�@~�7�ǋ����B?��9~ef��b�	T�H��Y;(Yf���N�{.$w���c������K�w�6��	��3���r��6�6�!Z�x0�ԍ�$~������!���"��ӑ����l��$��Ĥ�b��
|��"`�|%u�z�&:���{�f�Z�Q5��Q�T��)f��K/���"NW	�c�9vFЁ��ѣ��I�eF���?\��Pr�O����M^��liK�	�`���D�NN&1v�%7nt� a�����P,$��N5# �'DR%����I��]H�P�A��h�U����M�0��/Z�I��W%F���rS���ļCJ꩝�x��������Y�������o�����8���ת�1dܵ�lXz�o��Y����n
+\`5�$�WBtD���DV��� ���8>�L��mB�)g�a���oR�WI_���^'5���<jnʹ�$�{�hXc��������Fo��|M5�qQ2��٪��X�H�����M=�K�#}�H�4�o?+�?�C��~����fU+�Ϭ�W͖���(T*N�ᗄV%�⦘rі%�2��J�y����ş�����j��w1�A��x3q����Yzf�s��d�Ɨ+y��#LGx��}������E�)
�H�R&�>!��P�/w���e�#(U$J)�zɄXI���P���v���`ER��"L�ZY�f�P�v�����mM�'p�)7ip�S�=��!��
����C�b�x-ri��w�Ac\
s��iG�n���)��N���e��t�N�u(r��%#����,�O.,.�tV�?��_"�S*�����X6j�'�Z\�	9��FE�.�@���?�+�v�i�^ɠ*?�5�?j���h�YȪ6����|��߸�b+'4�0�v�eG��$�;GD.�ᇓ���8��[�����)��O"ы������m�
��Y��A�����%Ut��މ @��#,�_@eq�^�?n�o����:j����i=Z��H�$F��z���5��=s����鑭����&=�.���o�/�k{�H���Lc�2��s����I�и��
f�q�,��:�M�b����m�6���"�zS�2P�Qנ� ��n�NJ6�m4��*ѭ���"p�r͞dj�!.^��
��AR�;�aX�m��D�~��u��)�e�<f?�X�L�Sp9���J<��H���]ְX�j��7q����bȯ��"�{�}�컔Ez� &Ȉ�m�e�oC+b���ޢR�7����S�`^�x�1�9=k7I�كc��s_�A����A�D��ӕAQX�s����κQ��.�.���N�� J�΢�{��3/+ĳ�kL�MG�<{�����Jg���Gf|@�ͩ�� �\޷�$�,{?M��{��{���3����ԡ
�H���M��&������Q�~�P�Z�fh��d��;gG�f�(Kg��דI������m����� ����4st�ꨦF�QaђB����FZx��cױ��� �C���l;4�3�gG.E�ߐq��qP����+�GO�����D���Ԙ���~؂1����.eH��"����N~�6N�Z��sd^Na\QR_s)�����NȲ7��˿
�A�4��
�(��-疰����9��[[L�Уv�+K���q̨vր�0���4��/?ބ]�J��z��%�|�&� ����dhZ-H�ֿ@�4*���d�س7h���ct�?&�����Ӥ�2ϭ?��J�B�g{���� }��N�c����bÑC*���7mTU���lzDK$��x�k���}&s�xy�6A��)�BB���e�H���J��1���7�N�|��d�i}���4��Wm*=�E��-���:@����#����˲ޞ�P�(�x6ӁBY;���7V����Z�i��X�ؐ6���♟�5{Sc�bʎT����-�,���/n�ֹ #���o�8��oHv�3���(��œ�_.�z�룪��W&"�[X�fS#m_'�*��YW�8��O��S���3�b]xw8��
��d9���Ļ$���T	�6�����S�G*����.�Z��Yi�S-�؆�fd�#�G��:k���?*ɝ��D]��c:��`K�;��u�5]~ZZn�ޓ|�������y��հd������wӁB�^��+���n�FLX��V�|���:V�Bn�����kQ�p�F0��������$AQ�\��X�0��zl��h�`L`mz�-Q�Hv�r���8��Mة֜j���u�[}6�ծ4>O�p3z[�%g���,�|���C�|��z�Z"���[l+��3�-��x�����'T�J7���\�Z;�(J�n�>E�X��ͤ��\&�.��
:&�����7;f#����do��̟��C�G�hZ��'Ψ�_h�Y���˹�x�X�/���7�-��r��I#p[���Q�i���萓�b�q^0Z�` '3^��JQ��̄����f����C�7�rc
��]L[����E���.2�}N���͙��b3rXk!Ǆ�� ������&����5�7�%��J��5{�E�%b2���9NN*���q7>���(���`�*^�J­�f�����h�L)@4̂�O��f�p,0Wk��J�����rC�;�3ޗ:� m3D���*:��Q��()ƚ�ɳ�G�@�
*C�\�*�	����՜�	_&m�mIU�c)QR�k�W>ld�c���^foyYi�?;AF
v&�O^d���������ڙ�(���2�c�cp��&2�rVEѰ�I$pZ��T��)������Y��f|u?��#��x�\�<��1k�����r-7�4S�< ���b<yi�>��l�˶�f�v���P����9�K����fGP��_�,�=P��f3������V�+�rx������<��S&���;��fBVu���� d�pZf��/j�i/���о�W�qΐςZZ�td�'�n��B~�w^Q���}R~h���#�r!l����cA�
��ė��u���d��U쩳�X�i�&�j�)ng-_�ĵCM��@�o��I��ch22���t�؍'�,�t���4C���	�X�8��N�_Փ.`�.)[8*���e��Q�����/�3$+����c��C֍�Y��L�H��I���#���e��ӣ&Ia6D˫�)��#�c9R9��DFuhw��C�uc&�$=�������v�x�hp�&�����\���vtU<bd�x\gV
)J�}L�B�[I��j�����ӧ��ge�cYO��5y=o�"3��X�`}�����$*O+j}�.�Ct��� =څ@�\���LEh��������1�` s�$ ��Ts�B�P���x�n֖-FcX��j!YC�kh�>�j��4��`��K{��|���r�ҩ�9��#�Aێ�{N��h}�.�i~��2�T�U�`~� ��B�������S˴�DuӋj�B�͆D�&]��IN�y�{�9��Ɓ��nBtW�]6�XT@ymz'��Y���i�Hy��=�\�"q1�#9��G곳S�5|֛{�`��r�ʏ��7�9����F�w
���.�bX�3<!G�d�[��m��uA���9�?�-X��c��N�N�_J�F5ѧ#3J i�������շ8�%�
�T]}� /!#u�B��ܮN@Q��zBM{��dsA����ҩ�^�geAj��֚	���{�r��%��g[��|g�s������b�����o��+����尼g$���j.9�Xp��z��|D�	�q(nOftw ��G��}V����g����R��e ͋�E�z}*#4cӤO�+����`ID'�����r��}�6#��ȳ_"a ��G�{d��q4|����d�kr\�5^���'fH�|s��.�n��>
���?�j�՚Oc�t�	�hK���a�ٝ��o��(MBC�i¹�.?���bl��١��r*�M3|Bb`�����\O�/<��v#����x�R���O�Nr�X3�cLj���S�Y��b�,,�p�α���d�@���i��{A���|�.�<�l��~{�?�,�?$���@7�+8��o��H�������7�~qW�֞\,S�[�}ꗤ�`5���?9���3B�0�2��Y��v���#=�HB��#�N��q����q�i�>As3|��搴	�jʊ�����lM���/JUS;��5�^ܱ1��ݵ�w'M�^WL�,,bb�y6ف-�۫uӌ���tOɴ�ߺ+��T�q�*�0A���n)ˏ[l0�v�L;1W����Q���c�r^>�#'-^db���֗�2�,=��~�Tiq��TJW��&�f/��1����y�K=�d�}&9LeI&�ȍ���N��6骃��~xC��z���$�?��|	�5z^�-����^N����EL���(��z���?m�n�B"�i��cu����$�6o�iT�HobըÚ���C��t"��9�pڵ���_["���x�+�#�~��1�ђ�6|�X��`3��ֻ�:�5l�%L���Ѧ�Y4����� 9�3�5�2n�Z��^�����������
.���=IJ���h���}I�_U.�I5�6\N2b2��6.#-��t�eO^��>mX���:nI�(�Ub��"��M"Q�����ɁBaAF����{�e?�M3d������P��k`���n��>Wm��+rԕ��4$���i��.��J�O`~��f���!!��I4�Q*@���=;�;�0���P��,��n���%d#�(�y���!�6>g;dP�j�V�M��L>�7�F����]�U���6v�ym��	�ʒ�։�d0��/kT����f�3,cxRtptv��_Qp8A�.�tBrTݴ�)��r(��j!���}�4�>Z:��y�n�s���y&Yj����t�m!��Oo+=�H[�G�B �Ec�C�d*$�A�	���Gq�M��sp�G�{��v��A@�*<���.a4�\FK��^eG�x#��h�ͪ���UȠ�;/,W���{l]^��z�8�_0|E�Y*�|�� �~I�H�Ļ#�q�gۇ�2�x�	��cC�?����D���5D[��8���9�z��&�qJǰ�)�h�i�3���;�a��g?�����ɿ����χtC�O��ub@b��]�3���7WO�ǀ���,����۬��mZ�e}��;M�DO`�@���1o�����m��Z�Bt\ث�Qs�:GG�3��'kQ�@a���wܭc2��4�%t���EU&@cv��!�\z2s�:+�I/R���y��zU�`�ϵ�����X�e=rgmh��D�U�<�|����dC�`����I��!`���I�O�BKu�>�G5Hw0�W�*�7����d�)T�tJ�a��t����# Oz�
 �6��%ٞ^�J+�D�!�w��2�P"�7}�u�ǃ���5{+sM������a����C��'��-Yw�#i�A���:�Y��\b�I%0�Zpma�%w2ћɋFeX����������#ə�N�����-�&�6�U`-7�ߤ�G��]Sf9Т$	wG��2U�hU��@��W�?\�jֹ^S���o��6t�M�V�,����V�F��u�!E�!]fo�#��[�$��3���/�˫t^ߙ����-���r芦�������g6*���D��5m)���G�K�ԃ�8��Ja��"�`��������jc�(�}�V�'Bj,5�L���'�
x�*M���a�P�J�ʺ��gl��GY�/��J��3Y��p�L�c,Z�Y=6��.P����^��"��s ̑~bm���#��	�X"]϶z�5��h��{ u�|�aĮ���^J�Z�vY�{Hn��:mʌҨyv<]�n��~S�L��¨{ni}�N��6,�@-{��Ur���S�&��ϔ���i=�t�/���/�Dq��Ǘ#@�]���mX�����u� 9��moL�ؔ� �~��7�'#������I�'����ri�f�.��q����/���Ll�����"�b�EI��5˶ �����7����<3�ג����k��Xd� ���Y��)\߹]J��'/`\����+܍$�=�#�8$��n���%�)�/}Î�ni�`�W�N�0l��F�ȞDp���/��N��Y��#�ܷF�W{�}�W�s�Z>�b�Q���6" l�F�
�֣��eb�	[TpT'�Ӈ�`0��7M�{�2�B3]p?��ʚ��̂� �H���;N,k�<����΋�;4�9�ZI'��)� d�U��!�h�_H�#�G��s���V���,�UE� n1l\vM`� ��@~����s��J��wZ};�������=�:S����E�1`�N�b�{i@��t��>�F�ߊ
#�Oq'�-���^
ز���I�q�k��`����V���|�0Q��#��.y��&�IK�^l��5r��(i\}�jJ����+:0� ��29���HHx� !3�C��VѦǆ����6շ2
ɣ��9:��\�,n��6��<T=-��\0i��=Py��$ϡ��.��0���8��$�W]#fq������n0'���L��Q-<O�t�Ȇ�Z�[A��U�.���p�~�̖X� S�ۆf�F�{��Wv��bI���돞��;����y(�S���~�TѰu��0u�Ȗ8_WK���3��c<��Ae�^�j��kV�գ
=�"O�,H�|\���j��[�>|:���o}��(5A��J��H��fJХw���Q���&�K���yba��:�E�(�b�j�o�y:~����/ %�2���q�p��Q4�+]{���Veb�����]���l;Tnh����=���v�,'���;��x��<D�%�1�F#f�4:�ȥWb#��h����f���&M�ȇ2!������;�8��Ox;�{��]nf�4���j���IP���o�
��*~{d�?��Gp�۱z���h"�V�C��/"O/=mK�t:6A�S���׾Z?�����6z��V�L^��d�;�	^
[�cXQx�����z�`���'���:�F�:�%�� ��@Sh�[���J�溪Ӎ(��R��}G��MS�Uy�#etpC�ZX���E ��c���aGi�Pnm�j�lx�c����1��q�׳�*�	�*��[=ڬ�%]R�m1��.;$30�+".����c�H�E����5P���Ng�#U�s�������>�D������Нê�dM�W~����Hi�#�7	WYg�x�㎐L=��:���y[���a�s� m�����2V��Z0���o8�{G}��f�1]�<���b�E�]���P�!���z$�o�/#G�y�T��=�Q%��_D�v��U��	�:�?>�IKdW�C,��r��6I5}v�^F��hT�l��4?�q������S���0�W*{��)U?�F |0���$b�'�YW׭"����G��[�I��b �>fn'$��x)e#��Bٍ��ox~�-T*�����ـd�4����o������"o&����+�ٵ�c��1�чU�n��H0B� <�����`��ކOt���R��hk���ģG�x���U�ߦT�f�g��9�!V�,|S�x��b6�{��jU֥0�Z�5'ߌ"�}*���}H��,�P�c:���?���L��>�*f������ٞ�&J{&�P\�3Ir�yYKė�Ů�$���v���ل�᭿�)Y��b��tϺdl�{S���]%�2'd�*ѷf@5˿�	�FJ�l�\g@�����^޻Tv�Հ
м��44���b,$�\Ӏ��w>Khye��8������$Ҳ��)�-��4�|o.M��L��l�Z�fqg-`h�d�?D��sh��J��Z?���s*�4�#0���=~� J(��܆�A�篢��;��{j�� y$ ;t؊Y���b�p��YRҰ���n��dmt�|G^oL z���Ϩ�
�ES�M��]/UQ������Zb�)5���w�Lb���0�EjU���x�%�8j��=��3�C#^?%�&�6e��%���!�! &�&�-z�
��@Μ�k�ά �Q�4��)�.2v���f���][�{�J�U��j�����{�J5x[���w���t݀��������]�K�ѽ�Ӳn���\�+y� >B��e�l��
���o���zlm�ޝq������M����.�D�<܀�ٴ�/���f�?_ �^��k9�|����?��W���k[=:Kj��'#��K�\=��ڙ`.����-RMo?�����[����E��2W�kz����D���L�C �!4��&6�fW�=��$���T3΄��4i$Τ�V�z�6��roK5Y_�y�t{k���Ņ`}w��Β�:!���Kt��c6_��ӣʡ뎓��Q��v���y��ڌ��H�wy�V���b����P���if���]UAR�xCrm�
U���OڨN�
Z��U�C����x
�c}f�y�\}��7W���{ZLsb=a��n�1� p�]\�F��w�=j}�]�^~�Хh��i1�4�,���'�8��l�̰�$��0�,}�k��-�e�"�s_�xfz�BS�������Y��^-�P&3`+�U sM�-T?�$�0���{v:��nTVF��G�µ�pC��2��_���L}�V���~��-�v#��Η��������LD�5����X��z�w�W܉�xw�E��ʛ�(������-7�i�Mğg��hT�����j�7����\�?�^��"�==�N*&��% $�b�]'��_md0�*��I?,�<��XC	H�	,~��@:���e��6��TA��?�ϝ�_��~t��&y�IC�S�a�(����ҟ��|��Q��+���!�0�彥7�����r2��Z]��$�/���d��H'5 �y�r����AwV�sF����#�y�oeV��0���M�u����Z����=��!ʵ�a�D�zPI�!Y�j�������7׋�@1S^�̎���_]o����g�*t��n	�)K��ϴj�!�7>=�-���"��1F
����r9����5[�Y�R�/?�
�QPtJ��y����.@?�c�N.nkfh���N���+RgGSl�_ ��)Q�O����P⋬��9��x'VF��f!
"�AM�������E�J�����&ggf(��	�$4�o�zj�^��kN�&�税\�'z�PV��}�+gU-/|2g�b�p?�1;������zz��V�W��yNϰ�	d/j�|����%P���߰>8��4�����W�kkS$�n�p< �|��9�#:�?J!͢�ϒAz]�y�-����E�@�����N�4fc}�߿��x�9VY��<�p�o�Z8��{�� *��)��[4�M�i���1F�p��� >ѡ�Y�#|bo)���^�Y$.��A��D�ˢ��/x|�MѬ���w�=�R`��iʙ���*�����Q�_g?�B�o��Z ��:�_�Ew���b���9�󏩔CX��t EG�O`�qq;��Xq�d(LQ�� uc=�خ�c�3�5B$�(������X��e65��㿷���쫢g�lʢ�"��yl!�5�~E�F��jP�W���"iW�r�L��c���`���y��%H�1���e�~vpx@�_�	m�b<�����lx�plp�,YW*�A��D�}ǧ{��Ӄ�K���C}��%�=E.EMb���'���!���2Ƙ��u:�V�Ӣ�ܛ�i6���i崪��f��f�������I
)ѓvs2 ��������-G��R��g����ma��6{񟃨v�v�S
�*Oc/�Q����3���0}���C/�Wr?Q`<�RgG�!�\j8Vh_ے����φ�0����m�mm��O1�%��ûV�n�J�C&�bY�B�o�B��r� ݔ+5�F���ñ7g�Xzco��+eQ�`Ɣ�M�(r�|���_i��h)緥�+�ٞ���:ld�1�����,�jWN~�t<����$�h{QK�,�J���t$\A���t��h�\�9L��˿G�r�QK��Qa��1��
ؽ��#��Z���/(�$� 6SX<�fZ1�����v�ۥ�
K��yC�\�)*��O���>����0�x�2rn��d#�6�׼}�; �{�4�72��9t<h�5]+���u�-���^��BU�i�?��:X"=e�D�n�z��[>�:�l�%� �vJt�A,|/�`��F"���`.�����b�v=[��> ��WA��U;v�Ia	��P�Q�zq��?r]�R]V 3�ث�7��%�B���4��rc�f��o6?a�g��W)�8���dr���?};�d��ѭu�����_=��;:R�a���n�uA�����I�FH3�`���;�x��~�z-��*��Z�e��b��G:8��S
�okV���L����Z_� �����b���!��(3���� x�%v����6j)⿲F
�zsN8]f��������#0k���M�)�����/�Bt�Ճ�	"�;�*��H>�{'��=���[u��"T�)�~h�A���f�����,���3D��M;����p(e�c��/���`�ohz�r%��槿Q�T,Dau�>={�7aa�ג+�~�<�~��9Ԣ�n	�(D�#!H{��3Dx����껼������32�% �`ǨJ��Ǜ�I]�#£xg�k�	[Nh:����sQm�<�<~?�'?�� 4W�����@s���,;ݾ�#��=I��@���~�?�GP�%d��*��u��yi�P�)mahw�÷g3������������@rz���8)	ԙ��w
���8��H�o�uo��U⍪O��=��Ss�^�.�m��؅���y���Q��H�q��3�}4'<�L��a��@�����)Y�. 5Į_:��5ZQ��j�-� ��W��!ϠtN��;�n%[]^��&꼙*��{���D5ˏ#�+����[h[{I�K��/�d/��S��=�T�/��n(�|��GC�vs� -Aǘ�Z?�5ѡ8�m�o�+US��Q�D�MٲB��#!�K��bQ��������,��J��������:&�Y}��a�z�<�8[O��/��`�����9l�dϞ���B����}��ϷO&ŁGY"�^4th,G��j�g8��'��L(�s�m��1?��g����F�s��T�$0�5�(3ᴒ��:�GMg�N��D�bP!Fw����0r�s��p}�p�4�
�Y�B��J~a� �Oc��=dܗp�%.��m��t�Ƴ�(�̱�{
�NY��x� �(�$�ϙ%I%�r��+�Es����iz�9�׊R��M��u�h��.*�o��s�՞`r�c�X]��D�1�@�Ohiy�p� ᄃQ�:u�	@?�j����e�(^������9D��"G��ST������j�S9=����Fi���k[�!۞	�5�v2?il��M�ܖЭ)`v�`^�PQ./x�����@�y��?u,�-k�� %�|���KxQ�Ĭ��� ξr��a^T�0�Ͳ��4FY�ֹdg���u���� %���?�w#Z���q�;���F| ��e|�h�QV*��'����ǒʭ�V���?���|�o-F٦b9ʹ��5b�����>�M���F��x�o"S�W���7��ڻ�ˌy �J3�G4�<5���h"��C�3��LG�Ŧ�v�D}x�9s;[���_S�TP�V�D� �.��^�m��uz�{鎮lzAɡ~A�ؔZ.g8����T����Tg���r�N�@�8Z�C�vB�s�̆�{Y3�n"��
��
����l�H�k����v�����n���O)�-v�'̰M�(��+L�Tz�8f�^����-���.��#�
�C��8�R�I��80ݽ';��($39k�=��D��tA��v�ˬ31����J�؝p���ܫ�6��o�)��Ӎ�`c�:>�逩�����h��?�Acs*�^!a�lXRl�w9���
R�;�p6��/h#�V�u2=*f�T̿ X3o��F;�*׃�g=vɜ���&<+�[/2z��|�����f����Ӌ'���T���N3�����B�����������J�ȱ$�����G�X�hr��b�^t�/�9V�	O��@10!���^��6
��j���>��)�y��u��(���7 B�S1�b�m=q&�	�(֠.��='�c h�F�Ҫ��C%Hb������+b��2�w�awQ���|=��0@��j��Y�o���G�g�d�ͼ��;p(�tt)�����-B�2�f���7���smTT0�@ʵw�YV����^���*&�5T�yWU:EtK��/4fW��:3nN��)�D��V,�R��E�θ�7C�bX'����7*��e4s��kV�B&Q.6�=an�/��*�Ɯ���XL^H�jud�}d�ئ�e��r���"0�é^JChu'P5��4f�s��f���X��0z��BaW����4U5��qui�2�vb�A���Lb�=FE�OPĢ���2����2��	�|�,�������WW���kW�T������=�����d��q���G9��B�����{�\���E��H=���EN�y,(�$�d�� ;��2� {ҋ"~�mòI���P'V̢%<	4��ަ�a�Ç��ޚ!��dmZ	�d0�˰$M������Q��gtH���9��|ll0a#U�;Ef1e�c�c&H̀�05Z����_�.d��
��i p]�ά*L\7����&2��Pn��i��k��[m��ڙW�rXB�@���l0���X���"��G_�֓���w�n�Ѹ��e�&r��7�t`vA�iyJ(��!�Ē�/��#��]��xu-a/��o�޽Ӽ|��E�����F\/r���"ߨ�f�9�t,�W�0��I�N��4�A_v�x���
�h})�nWW��q�UH��R���ƒ׾�@{���G��;$����qO�'��b}�Y]'�R�x�u�w �͖ /��,7D����r�V�R���
��Mȏ�x;1@���ibZҁ=k���֐�3
-'j��f�*D��
ӷY�����!4�K���Qu��u�uo��ٮ
���Eh�L���vI��Y:	~e:���w�r�i�Xѯk1/V���#��ʎ����Ƭ�;��r����˃]��m�bTB,�!0mIu��݌E��̳�٥�������̷�6����:����3#F��PM9��,��a��m��"LT�d���;�&� 0�F�����ѥ�w%!��35<��^��%��m�}��5/�����5��5�@�\����!a-�s�,���C�z%9��d_���u�7��n��h�@�9�L���	CX諓�&oZM�;z6 t��
��{q�߂o�: E{-�Jz5��׿�R��YhHl�F	Ðh��*�͑��4fu=�'���~2po�WOj��.��u��.�,-d1y����
�U��K�!n�B?tM��U0���}(�����q�pf?"��],]s��$.��! ���[��,s7�9�rpm(*���4V%U�۬B�L��W��اJz{�tC�q��5��ذaY�g�٥C�a(/�G� ��x�b�z�F���b+�X����-�\)�}�CO��B@�Kÿ6?�*Uw[����0�#c#9c5��C���Y�|t��!���Ӱ���Kŝ���$"��(�~�^KJ�k�i+��>��KJ����I�{����lo�x<߅�u�9j�P��/�`�� XJo9j~�Z1כ�@]$֒Я����p��U�!h@s"e1���p&P(��ѡ��[q>���-��;;�|𬄿O���� J���q���9_��R�!�Ԩ���8�T��	6��}���%ދ*������̶�L�y��pI������ �A6�΀�:�}w���a'�fd��YJ�l�Kdk�rP[#��"ell��lخ�v�H��q�-ꩭ��Q� PZ�s<�'����Ӡv�4an�_5��O���(ց��~��岹re=}j�?V�w�::X��tZ���~y���
¹c��m����3X��=3�^�|M�N��g/�/;�s�B0'>=�1��qq��Q�q�^y������T�5|s���r' 2���ncA{Mڣ)K�,���k �{4�	p�I�ov��p���~�T������}c���=��A����1q�ӕ�6K��
�U3��,��ؼ��wn� 1�P�r�}[Xw�%e�����!�ֿ�7%K4_�]�?ܽ�F��h~2����1��J4Q�9��"��e�G0�(��.O}��]�oU�qn�.7����]��l��;�����N�7-��B��3b����ޥ�|�@N�J:������)r;S��k�����+a��jX}��>�s��H��#t�Q]��D��S������:`�W�X>�,�W�ڶ�6�4�\Y}�&�6�y�o�N�ZA��"�~A�����9�|���%�@+���;3G�a����lx4k��S��;OzFN<;~��&���z��m��׃_IG��9J��-Ag\l6�$}Y̰�Ï���j��_�ч�B�nk����kY�0�K?5\Q�������M�Ւ5L���*շ�q��*�wW���N�)�Z�}���C}Ck1�>]Զ\����]#�^�8=�@����ڰfX���jcgP@���o����9�[\�-�e���R���1��0M>��W��^K���vߏA���>S�R.v<,�_���3��J���=2�2m�B��������*�
%Ԁ�:������_D�[�l��� ��bÅ9�����c��𑱇u_
kD�ea��|zʅui�h`�S$�D��K V)}Zhz����8G���y��L	#J��{2���T�hN��i[�����Z���Ph�w����E컿�)8t�n�h�w�D��zM���U.��׋�c,,4����Xau�/���z���Ȥ؂�:�:�<�с�lQ�p�����v��wglM�+>Z��A�O�s��y�z�'IR����*J��]�B(�����Y�+�s �Hb4���/�Ѱh��(�0��A�!6.!����%!���!�`�7>Y��v�e���-e� �!MIx$sK���L����X�)��V���g�H@�z����m�~��F<_C1��@݇�����YY��=�'pr=9ӊm���:"]�$r��qG�$I�۹������Y@#�+P���Ӑ� ����ƌ���@��n��F.���Hrm�rc)��c��A?@�:J\9;��i�0�ʧ��2e[�n����j�Ê�����g!�O�[4�_�oj7�ܺ&�������
^��>��tsرgs4?�v��z�7머�	6�^�O�� 6�܃��6���d�b*�I佯Rӆ9N�u�i)�xG�{�Q�
����XV?E�7k������"�딖���V�i�;^%��v�$����F��}�A2��]��ȟ�� Ô~`���B�.p�p3�����(S��3\��9�F���;��ᣠ`�QoUT�e����;u�w;0x!c5� �����)0�D��_�=w���zb�->z�(SF�j�{�r��y��琫��mpy:�Z�7�S�2��������̽��,ݭoV-�<R��B�D�]j�,�莬ޑɅ��Ԙ���P(�
P9JJ�!�s
5����u��M�X�*���5>�Qyғ�F�<�n�!%͝�<P��V"TW(�Z-:b����v0&�B��t�'����\i�iU��i<O <y�ןU�(_�j+_^�=>����TҺ�)#/_�D����:���|i��w�b�*o�ĵ���W��(�"�E��֍^��p���iV�ۢ1��(��KA��db����]�^5��k7��&���zC��r}Ci#fe�>���� ^�L�5�a>��@��G��jV2��ڎ�Jp7�A����>�^��'=Dώc+�0~O�QF*ya���k�F������G�������j?�w(�_�%��yD��ʮ�����i��^h=���C�>�q�1R�h? �S�ϤJ��_�6J���ki��wkl�I��|7*��H�������H�C��P�Ր�|\�Ԡº����0L�Ja,H?�� 7�����U���Q�˷������,(^> �Nizz231�ت�^|��1viQ����M�ᵰ/R��6�7�F�ms�u�u����Jr��'A��g��r̾�oCc�Q��}�2�u�S��gy�i�" ����*Hn&��ju�!:���B�?�; /G8����$�X}L?�6��~�W�*I��i�Y����m&q���J�}9�*Q�<�����}ؙ�������D�zҁ{X�Wb���>�\��\Ii����_����"�\�J��2V=�欈�ܠ��b��FQ�ƀ7fb�~.�[�(p;- �{p����k#�&���8���;tJ�Y�&$^i?nt��m5Ǫ���+�]�O"��,Q��+`yй6�8"�=��;�@g��;�:#;�C����k]��fJif��f�)"55,�)C��`�9�я���l�%a���5������ ��\���,{A�!=˷���(�\���-V�tM��*�=�T��xʢ��w�s��Y��7Pp�����_=a�a�R�z���]���o�6��>}�B�tW��-P�M����W����1�<��Ip�����MLWi�i��
��Xܠ����Y#�;��S~�_/Ñ[.4�Y]qj�-g����`;/~�r��32И�B���6�'��v�v1!}����Km�q��t2Jq��b�~YiP�n��Z,^��uq䑓�?�U4?���|6-s�z���WJ�>fs-�k�K`��DW'����g<򃭝��������DKG-��r�gx��(�V��%����6�ԝ ���8)x��
|Q�K
��t�/1�|�~���������{��@�q�-TD�(e���ݽ�j��`r'�w�k��ъC�؟2~t�Ou�oU�p9�-D��~+����m9��'�kZ��5���=�H����ŕ�#��GsWf���3+�;&�/�=��yw��gr|'���������NP(�.?3�0ř!�+P��%�@��+DD?���g�H���g
��$�`���zM���ȍ���MfN�pO�7S��n/gZ��z1%�|d6S��~GzqH�7�I�t%y����o	mگ`pӥ�����;����E�ાx�;˰�����C��أ�alV���,��8�K��G�0ɜuZD:8�⚔*T�N.��%1-rZ+�n�2�ΰ�����~���m��'.6����������L:|J��;*��.9a<�����Sq�I�JA2��#~�*�O�3��M��|ӹ�-�y�qFab�hҿƗ/�� ��F&0�l��@o!b�
-���1��㠛~��j|�	�<����?Z���;���Qc�N(k�U�O
���D�٘��ԛ��H��nh2Y�6��M���n֊��N�������ova���\<4���>q-Ò��5�+{�ppk(�#Gk��b���_W�d��A�W����������ߑ̈�]ON.���	��{q���T��8��tIAW�������	���m6��Qz�dS[ɬЏ0CG.�4��I��loH�|N��4�3��ȥ�� �W��'�5����-'���Q�KZ�Q�0>�b%��*����Bi^�t	&/RJz��e�BA)6��h<�"�$�l�,����W1�=�#��l?o���O�q�=�r�[���p�w�D�H/������DX���C� ���8��c�㺊=��4��
�6#���,[O�c�k��lTb3 �̶�F�ml�Lc�1��n�zR�A;�*6ƶ��[�&�b���㟘��ޏ�bg0,C�u�tr�ݭ���Ʉ�n(��@N�U��';&xѠs�*M���.�i��a�&�c�f{�sG�em��vq�eU�W��z`Uj:�z���n�,�noe�q���&�/ޟ���3s����VڼZ�!�yc�t�b�bb�$�J��=q8������i�G���I��1���h�v���|=���XY�j;�I�8�m���f��Z���p:'��^Fk��C����om�4If��e�c�\���R�x�Kr�}�|+����t��1a�\�sb8�FY'*.�/%��t�"�y��6ga��T^|�pY�c�]"ȏ\ϓ��@�j��Hk�����r'�M7zQu�}�,^��������0�F{W����]^�s�oˑ�x��:r�Y�2s�t�[C�d�IK
<%(;��M>Ԭf~nf�.�XC�'�C���GJ�ɊG�����t����щ�٭�~B�,^,��%�R4�%���/��S!��+83��j�D+}k�H�?��A4�B�/��>mq�>`�lG�w�yI�%��!�k}��t�;����ܨ�&���:3:y�A5�a��$�o,7���x��t�kG���a_�џ�3�a8������eRB����.�A���@M���L[f�ۇa��kk��0���>�����]!-�	��՝77y�o�t:�
͢1��+���B[.�^jԫN<���.�� �����OX��'CI�u��ζ�9�k��T)�i�j⪼�;D���w#���̮A+����X�AxqɜQN���W�fp�����ؤl�D
>�e!4q�1�� �cS����jL���E7YAe��:�Þ��	K�G"�f�K��a��j��17�f$4�뱰'3*�c=A�mL=�t����܆�E�� [vhE�y�u���`��aU�7���ڭ��S��l.%�w��ګ����R�,�.����z��ZkTf���=��J�=��T�9l��[F�+�� :D��oe�L�B��+P��ܻ�����R4�\���?O[?��&�S�����S{h�\/�ډh��R�Tq�O��\G"��:2q�ȱۑU}]�:t��
D��,��D�m�q[ÿ�����E�!��a�ě�H�lTa����Y�d�w�RM��;�tPN�B�I���4�C��(�Ŏ;��i\¨�޷��1jCo�K��ȔN��:��m�T�Ug�Mf�0\�DR)}���>��%\:r��fo����|Iy�,��`�"��Z���|�޴cjp�:�"��L]�@ȮY�Y�����~\�w�tY�я֍�� ��)����j��+̣m���!Ў���V��$y��lxB��2�s�f@¾~[�x5�^9�Г�p�� �z�!1�۾r'-BL4����C���#@�F3�!���6��^���g�:?�L$��5��Bf�It0mS�ZF�ŀ��=��U�ט���0��s����G�qO�B �{9��:j����ۨ"�i��,�����+�X?������S�&�\ଏZ�����p"����s@���r<� �M�� ��u�ᩩ~�<(;s3^�-zOaR�UQ8�����FyD��B��ߢl��IA�J�p���s�\���K�C��Qع�B�	Y`�p$iMC$�M�I�;�}�Fu���]�y&�R9�h�^P���Vm:K���x�,������������"-��'�vhG�1�\�o��k�4c����J#jf�k�KM�J�� r���	s@���u�](�6U��m��G7�0��n۫^�ѳ�o��̆������5J�(��SM�Wr�Y�P�d�	�b�C��K'0t�c��⇋�m�*&���ki�IhS}Ɵ��C �v�D�)����)$�t�r7=.�7�W3+-�U'˅�+��\^�F"jN��8p/-P0�~X��ʤ��49��H��V#�v� ��"3X��������R��hHM5~��jy	I|S�(���˻�\B� �mZ�PM|A��nP7�+8�#�
�y�C�"�[JH�oGX�!�[>Z@n����l��I�@�y����!m�>�Z�W���o����G �_q�Nj�2���$!g���L�Ǘ��G����O��H��/P໸����b���Z%HR.��9#k�E
5�:����D���4�s��3~�6�C��U^����DU,{��4�9�0t�Q�^�Z:�;��3����e�
plCRjՠ!D��������-��*�M\��l�X�<��ە�uێzd� �^[�% �(l�'�](+�pEǒD�-K(:�:�w}�Л�w�@�,�Ert{�a�ś�f9�#
;��#ׄ�e����aA�q�;����1'q��-���9�:��fC��E��!��ф�@��KϜe���ǵ�:tI��@�h3\�X�X{�Ky��Z�l+�EC!�17k׊MX�v�w���:HҒ��3?�0'��4���?zz��Y�f`���v�2�W�iz�cI��X���5jF�LI��+�F�?�T��{G��`�і�v�����������n�4ĸ���o�<)ɽ���ږEpP�VKa4��M�y��	=�A��s�,@<u�$�����a�0���*��@�O��U},	1�Grh�s�j���k� ńd�ڪ�Ɋ!I��z��5��!ni5*��:�M��MV�ۻk��ۄ�<�~c?�ݔ}��ߺ6�$���5�ۀ�ܙ�:�F)���b}�C$��p�()fCqY|20������-�f�s�Bɽ$�+wvϡ} ��M�J��$��xvP'���.򤙡g'���X�} ^m�n��)Ys�b!+�ڧ bQ3{�������]p$k�S��9c�M~�`##Ӄ���*�8p�3e�E������U��Ɯ�!2�u�n�b�w�������j��s�,�'���1��
q,��8��� )���w�'��܉�??�MB�֧U*��U�P��6C6hn���~�����/��e?'�I�i3����];��<kIa�����/7�[r�S��s6yj�qqLP�,ȉ�$pv$��xʞ	l�@�z������¢1v(.IgNd�l7P���仆�Yvwzx���b\d5�����{0����ė�����{(!� �I~e÷O9v�e(~��m��w��M��6�e�T�D�e�-s��ɴjB��m]���r�� x�+Z�?�8|��_�dVT6�_� ��fE�����9o��H��{�%�u���9����R���Urq�ؓ��)��#��b&N#��<	&]k��^ G���,F�c�j�)!�X��J��=(���yB�[���rr�w#�a��X}�ٰ�6��zH��ū��+y(��S2`6۪N��'H�mU�Pw�>����H����ݑ�_���O�c��=��)�G��� �#��Hd1��5���-�a=.�`����<5a�^���n>�7�ԹN��Wn�D������]���,�>�4�E��)su{���٬a��Nb���L�Ͷ Q<:��cZy9�zu�.&z��b =Z�Zus�L�8.�56|��i�#D�0;�쾂�;qE����|��K������>�A�f�3�t��R�Y��S�J/��K~L��ga (QxY����7а���j �07;sHIYQE�ޣ$:tI�+�4��ɢ�tQҤ
cKlz�
��')�m���[Ԝ��ؘ�'�l�L�αr�ف�U����������B�ħ��K����#�k�-�@�D����b��g��Mw� ��ԁ	��oiu�oi�Y^u��Tl#�Q�� ���"�@����u��FE^�H�(رDp��n�p�L�ί2�YNw��w@ei�Y7T z��by2��m�m0��DRc��q�7���;x4l�(�zr2��VU/\|X��&ᨄ{������D��ɰcF���.�`�}�b2�W`���Զ���$�����L�����DS�t����>˟�dq�+[��.��׺5g}��>�6qTQ�E�7��dr0ǰ�ޛ�C���x8⺒o����B΄Љ�zz�"7�����g�'@po�F˻�I�c��Wr}�]��[�C<Ӛ�=iR���8�#����Ub@*yq�1dmuH�P/��!�F
+BFAA�eoYy:�&�q��OX�����F�Ŗ�?�+�i��O�4VU�,�-������i�,%7�҆#��Z_]�-SW8�wc���X��\O�<��棗��>J�C~����;O4Gw����uH�ߍ��� �[�m�-re �4P7�ɒBr���8/��A�=Hm�Zh_9j���m=�T�m}	�ڔ}hP��8���A�i2h�=Ӆd<����&V�'X���o����O�%�퍋� ��5t�h�^���NB��գ��#k^a��,o�X]#kOuI��X�;z�*��&�=�G7ť�P������V}��;�֮o e�@E�.�m��w���u�0����Z�i��loSx��v��l�#��[�͌i�ysx�)�Cϝ7\�Nt�jK���_�{�؂��"V/�߱����k���R 3b~r�N<t�!ר��I�Zrr$AP����X��@����,���k���Fe*6yh�W�c�ĩE��K���dg�޽�DUA�ρauǬ�T���q���u ����D�|9� �gIM����5���n��+:�u�� cX(:�:3��a��o2��ñw+�AH�) �c��:]G����iy�e6S_xdr&�Xۣ�7�h�����7l�rv��7����mkw�°U"���lq�׿:tf�c���z�t���};�'��4���Ԁamp�;&�9Տ�x��;e7�����eX�طz��ya<9%�qjaa�F�GtGⓜ݊U�a)��LF��G����׭ܻ�&U��pOF�g._z�T����Զ���V=�|%·��e�?|6��u�e�7p���'k�)�l��J�@J_0q����I��n��=���TRc)a�I�A�[��{3��y6<F�e����f�IAf;��L^���%�2OibQͶ�[�';����]\3�j�������<O$��D�z�_�)�nL5�Ì ���fŰ��xUx�p	�Rj}�K�PI7_��i.	!��Sf���b�*����v�x#o*WR�n�<I�����L>ɬ�Hn�ձ��N�1.��'�\��ݐ8���"��\l"�t�k0�UQ	8ki���)��d�q�����ߴ���Bm #�e\�+I�X��GQ���9X���b�u��ߋ�Xl:1����v�@�'Nt��j��ɍ�Y�7��5�Y�o�Q����%�㽍��Î�_�c��-���"a��ck*���Ȫ�Η���iʂ@��V��d�ױ*"pR��R���B��L��R�!]�(ܳ��m��.�Ŏ���E�$˂vx�v�����HX�H��:w� ����ې���D�oZ2k%��e�u�h&�q�b�k����x�?�vs3I1^�xs\�.xW���
��$^˅̶+>'�!�	 ̒�R��,/�dX1{�J��O�~y`�nw�p+�IGp����ZtyJ��΄w�D���-Zܔ�1+�5��8H|�ѩd<��>��Pv���9�y�`{=����)=W'�RW�E�Q���Iw�N	��JCB>Pk�����#+������k^���WD��D��Y3+&����Ǿ�7��ڮ
��U>"�z�z�t|�h��]v'�RO�k3��j�X�ΰT̰�dof��D����ᰛ��&�r-����ڰ�-������kl>^H�h=?H	�(h��=�����B���C	��� ���H�A5\H����г�fW} ��`���1�:��J��=�Z��ʾM1��My��9.�"Y�s�s�������2�4�����Y,��-��qM)|�+�W�;�U�UG��D�ʥ�%�0_�.D���nF&�Jٝ�[@o҅44N����u����=��V��E3�q
4
���B�=@ևjpRc6��1^$�R]����.�C��zS���z�3�kh�ZQ�6�k]koԳ9��hC*r2�������5�<���ܓ=q��<���|Hޡl�{TA�r�Y2N�5����)lz5� ��ڴ��W���׆gN[2~�G1�@1���`U�b�Fӗ�'�M�`�9|޽�ζ���`����9ST��H �c��fR-\pT�KzD%�x�2|dF���5�ؗ=t pޥ=|_(�/����nP��V��:��7o����&��k�b�T��-�{�U#��>�����=�K6<�NpuS6��/&�ak�\:x��fe΀`p�ɛ�$����|��y��(މGMT���G)p@5�#��b����B4�'��O�st�h��)v^ X�'�)'�%x��6��T�A��u9�,�$�I�K�M�����l���ĀkG�o\�H۝^#g*������	�#Ѥ
����w|;�>7�q@$�J�Y���Ϋ๢�4�tw��[$�4�	�Km���ң�tzr�J�a��
gb�;sð�c����m0�SV�� w����Wז�Ų����C�u�Ph��y[�+�GZK��	��8n{*�۸\&Y��:R@O�M�������i�K�20��C���鞱���j-���3,t���k�6�+TQ�S��x�]���!�>"�߬
Zԓ�c�͆�N�Z�Y[M��]���u-,J�����B8B.z1	�Q}O)��|qtl6@=�����GO�,@��� ��\M��l�0�n��X �5�/}և=U���Zw8�o�B��yY�u�+m���#����l'���Wg��q�0 d�������$g����h�AR��w5��yG����!!����C¤�qNĺ3��8qmT��3�Vvzy�T���^�p����~>�C_THc���w�(F�U_��Ib�mzcr�tC�DX��3X!;�]�n����`��0��y�*z��%70����;�%��\7��X���!�g����`�Ok�hʹ���◪Ŀ	��P�1CU���~>P��������5=u!(�h�H�`��|�l8ʞ�{4��D np�y�ñ�>�tX������qL�pj�e�M��sPoP2\�Ɣ#���&nۚ֕z�F	'}C!��`>��725^z�qTu��DG����Q��Aj�SR��;�+��7���ŧ����*a&���B�����)�xcsk(��+gtj�n����stG��=b�7O��
���b[P���T� ���|E��羁H4g)�Hpc�p�4�����-:�sL�G��X�F���6)��qcIF��l�
��WD`S 5�\ӹ�kk7BD��?���"�	�#1˓t��`PsY#�7�l_�w��^�Q�_�A�>L�Ho���Y��np.i��v�$��U@p�V3�Ħ9/�hV�G�X��?��c�(�J�кVn�`K���������;װ���[r<_�v���CLV�iqY�Q���t���SZ5�3Lr�^@/W;~�C�?��2��-�u�}��^�[�L���4���l��'2�8�!yX}������^��SL�;5���N�����¾|ɱ�a֐��4t�l�����
��y��B��U ��ל��%�Y=�tr�m��V�U�(z���E�e�Y�z����fĨ�����m7]���
�0�}:�M��r��m�q;��<�@�~�e�5R����?>�aO`�>�z(~i
��␒�F��#ܹhc�6Ï��fz҉Y̫,�h������K�ىN;�*R'�Κ>b��F5���Ke�~��]� ��Xw��/9�Q?M��9�����*%�J/�O��n�� FG�W_pE����i�#߿ν��+ ����[n��� �[%�籕���@�)�ʭ�ߍ7�iR[�Bľ����(R�վ+b2P�!(d_�t�v�v�����������߼��n3��;�P����C�o ��é����
������k����V��jh��� �Q
�1>#��F�����KUD��ܷbB~C�z�6����Z��y���U����z��^���us����_�
�Oƛ@b���i������L}L���x���9�+��\�s=ƪE���u�Z��4o�EV�`��m1�]�d�UQ�Ϧ,��q�i��o�A�R}���-p�vU*&��FF��zW��u��!S�~bc��y�%�;&?a���bz�Ί(E=4JnS}�j���=
��[���K"!û_ ",�(�>w0����`��H����r�|�6�M ��G��J��W-�a2s8X����qr,F��C��H/�j8q��}�ͣ5���V��8�}m�����u�i~�v@ɟ>oQ%/G��KW1�`���4��Ys����NsC�#�^�F?�t�H����!�j��g��V\����7�'A	L�۲��AV��5���5A�S0�����9ȫ}����-�r��`L"ln1}[�5�G�թv~捎,�V�$a��S�_1�y���0�xF��r�s&��B��-������Fp���Q���9�
�?����xF%�'�1Z���̛fX�7��E�x�-��؟�+Ku,�BHܮ$O��TҰ�g�=�>��t)m�~o-��+�����U:��nX�,ԩ�	DD��_PHA���ĆSoa����l���g"��\�zR��nt�<cꚠf�u�IaI���I$(���92˽w7�TB�ȶ�H:��
+��E�U�4 d0����3�t*Q�&7��ZL"�,sM,�٨v���"��GV�G�9�~�<����57>NF������t��A�z#�L{��>�����o<ޘ���B�,.H�_P�n4O)�ji�9D_]N�86w�'d�~��ǏͲ�O�&,��?�z��F촏�Uq:���P���h�'{ж��H)\�+����,��F��ZXA����_\�a�G�N ]6��0:�UX�P�>F5�x�LB� H�B��ԤC���a�ޞ�e�s���?d�us}5c��zr��'�[�V�y�s�Y�]��6ʤu��T��L�2;��|~7J�v.!����d�Z�(��Lm�b�n���G�x��/"׃�D���F�B�#^U��nč�.5�LN�ȍ-���%�@��i�=�=3��9���9����U��`R��\+�P��}P�r��d�a:L~��Y����`��5+{VQ(0L�Ca��qn���d�ɴ��5^`���q����Ԟ���2��b^@�-���$���������e�A��և_G�l9jf{�+�����w�� {i�}n��� y?g�^��|N��+����$q�E54�aA�O��Y�ɵ��+�*����ޟM=܏�YvO�P��R�[�$I�\x>^J��N��)Eؑ³چ*�|�<��Sk�!���rD�j���_��c���	~MIn�WD�HM� �7$Z8)WA�|���%$����_P�qgmo��,͚�I�Q�J�*���$��J���6���̩��
��3Ǣ&i�`�FT8#y��Yh��x;��`[E�G9�*���`�͙S�C_�Hm�po:�[�(�u@e�����R`@.�If`G&Cȭ���'�x����'���L���M�Y�CXKs6���)���}�ad<E�հ�X�/O(������>5�u|xEv L�֚�
�XŠi���A!�2�G��*��lN��D@����3e��4&)m�!n=s#b��S�D�����=�Wg�4�����P���\�K�3��\�4�?�k��-��2c���<z��ϧ�����0 �Җ��E4� �y���9�� Pϋ���O��:�UH՞�Ѽ�6���Z�;�V��̟W�ӣ���E
(���$��9gв���ЊX⧋�7&�����vK��,B���jj�~&AP�5��>��f{B�b�>������]�o�q��]��J���X:�$V�,��e|�����O9��̋��������q��O4[�b��}0˪w�Ո)=���@t����/���
Jt�6�?���C)i�R����Gb�� 7m�B(��E~u���4TIgu�`�a#.��I�Ȗ�ļ��@=B4�m�E�?��o;��&��[a~r�
���q�ir�q�G�s��e�J4_�/�P��	��=�͕o~�K�]g�c�">�hm��mu�3�-��r�闎��T6A���Ɩ�*sF	�w�.b'�`���i}�@�hL�U;�%�vQ��l��vv�)��vk�ǡ�$#	����k,z�E�՝\�k�;�`�_��#Mq����3�@��/�CN7G
�t�`�J���I����W��������<'pX�E͎��b�&����C$��O�̎rm�8Y��r���<������̘	�}��TF�ӑ���qK٣(���G~��������OL��E�َL��֦�F04l�Ep�b~aS3�4�� W:�c��6���W=fpm��|[y�nw4�֒9��z�S��e��s6[��=�(7R�{iUA��n�Lz@�U�$�j�JXUu�Pt����6w�Y���H�q���������ϲ���xq�W�T����vnPmӐ��#C�3��^���c<���i�9 �K��*6c.M$�H*�vm�?+ve�#W�w[y��"��۾����s9�i�6���ޗ ʝ�8���B��Yl�,V�'[bmR��V�7\�2��v�2���|�ME�rIS��L��4�>�(�@��v��5��.��O�'��2�^lw��F[�+��G�C��8$�Wc�/5���^ ･�M$���_��;��jW��]دm��C04�@a]lF]����xt�S:%��h!�O�5}�ˠ��S���{N0��q���#&�3p�;���3Zw:s0�XhK�ZHTz�Vw9�]�>4�*\~@>P�h�r>�׌�ݣ���N��S��ۓ����n��dPC>���#�C�Vy$p�t��ja�!���O�w*M�k��X��<`Kk%�� �0��|�p�|t۶��ƕaii�2n���=�A�зyB)��M�H4�i}���9��&\��]�|�ٺ�M��xP�8�2:��� ���7(�X�R9yՕP��~����3�sC�b�w�K^}p^�=�o��DiM��ds ěCm�0�=���аS���̱�}�E�M8���hL��3E�*=^�#�*��"��s�c.�v�z�{�$���m�b{;��P��$<D�X�=&�l���� �&��2|b|z����7��t��z&P1��Rf�|H��74��b\R�.=Dߵ��#��@�u1{\0��:�g�}�/��&�b��߀!����.���X�� m��JC+�.)��J�t�|��2��Y�0�.��ga�`�:�t-{�'��ދ�$s�"�3�
����Be��29����R��i\�b� s$�1V
h�]���8݈���{[�{����eڴ	~�V�%��׈L
��sJ�ζJ���Y��J�����* ӵ�ԗ$����K\~�E���\f�(��AI�V���8�0�j������=�7���B6�d�"�n�c���8���t��m�E�r6~���I�o���@*.�B���f����噮�3B�1Cv��ʁ7��x�߄o�s��$�-�ߦ���]�Z������ջ̇�nK^�����F,wE(��*����N3���>�>
o�1'>ϡ�P a�F��TO����@S�̕MZK�m���H��vAH��@	̒$���h|!p���]��d��9�>��^I~�?D�K�;�/���_���S�mH兛�_��e�������h�E��DI���rC�ۗK�Z����Hr���u��1�#�]@�j|���dOW�\@�y�6 :��;�H�i|�r"�Ɗa�~9����4����-&T<vc��̩Ӛkla箁�/�)��UdG��H&?�V�ԺsYq���)S�s��]�
��D:艡�H���&��u��!�� 5�˸�BGu�k���oqh�[l�x6t�'��V+ث�"N/��@��i�EL@�9�V���5�ӗ+��sH�pdrzZ�[�k�)j����L��*����>��aL������=%�c�I�9���&/}^�������]�|u�x)I�3��P'|��{�GvP���zb��U��Q7�pe{�C:-�2�^�R�J�m}���s`=`��p2�eS}�<���k���[���f[IQ��Aw��kx]�nq�k�b&��?��)���<�9�*E�XYQ��|@��8�&�-H����<β��P�k���'*����U�,C�L$z�����EazX�?�6.���=,�=��8i�Y�?�Y"��;�W ���}P	\o��~;������t6�ƤsE��y����� LO�J���1)����~W\�Y��P
�o!��ǃec]�_ꧥ,o`���
�����
�x���Ub�Z^n<�kg�	7G�s�P;mi�ަϪ��e��f�|!����\��U\>̙i���!��CX�Y10�������M��^��^o�B`f ��Vp�f��"�y/T���;5_��p+�*z�}���/s�^4����R�m��v��O�1=��@M����"ϧ`�C�ߤ��p������@�qB�C%F�ܴ�@�8H�]I�ʼ���ZM�!�K�c��F���yϬ�>��o�ǚ�a�̷��]/R�����	���.E�:#.8j�_7��\�p]��f|�_��{\�3+�o}~[����k����:�c����{%������Q�Z��|ϯ�<��Jp�����ja�\)�a�b�
q6;Ō�����{�^A�tu���	��&��Ŀ6"��0�� +�lX\�Tg�^{*YyT�J*��u��e�L���k� �����];ӡ�e�%3�����S�щ6B�����������z����h%��י��HB�kZ����@�_��=B����%��t	<���
��͓xW��r�h��|ʷp;'@��u�~�Tmtyn��� ����\�0�V0 w��v_�xZ���|e�[�-�:�K)"M�s���+��YѨ��8��M<U���L��;�� W�B5�r��1�A
,�)m�L_В�UŸ���d�{��ة`_���otg�t�y{��X�W~9��Ɓ��k��i�ʟ�J��!9ߧ���-/�9?�΂1A�t������/�'�|�dJh�'e������ǹ��kK5^������@����'�-��YhYޞ�S�F�:�2 ���� �-����� ނs�;W�l�p$�� ��&}��!D�_j�0�gi��l5�F*���m��d�H`M��iݪp�4<g�0R��� ��#-&�k��K��]��/�/=@*7���IS8�Gm�w��~]�Uc�o&��(����j�ЪJ%g�V�#7��Y��E?⻌���ű���;>S	����7��b���c�<���Z����d��� Ip�,�����f�Jv;S�����y"�S��b�~3��>�IZ;�>#��~้Z�Wcmeia�z��pW�]�d��c����)�EhعH��Q𐡼��#��䗕���mႲJ�BeM#��h�f�xT'.�6=�Fd��!n`�&n
_�љ�a��W���zK��.a���:;`�)�S"!�+�B�=�؃�z*��`τ[m��	�6�ځ�#B�xYg�ar��H��ȁO��4wD^�r�q���<�W�;1"�×�{$#�^o@��{�Fi�ɤ͟�[4S�N�S����t��=���ɺr�m�`��7���檤P�F]P'�Ȁz
���`g�#����jP!�6�����a���";��/����x����}�΂W�@�s>f
�oL9)�K�h��gJlG�gu���xD�/��;�邟�ڄϸ���G7i���M��T������ D�s�-
(N05��ݦ�x���8�Q��o�C#2B�.J��c�[ @#�$<�9�\�
��gf�J�)�){���@�$�t�s@�����K-k�{�A>��~�� m.n�1�.�YƦ�cf4@ ^�S�O *w��{��h�����P�9�ğ�ֹu�.Ϳ�����w3I���:��R~�|2���J�R,ԱZ74R��3A�v�Xt�ʓ�ꔔ� d�����a!�44ACuV������{�,�[��?�^�)ѫ����?��{���`���2�m���;.��T<bDui�(&� ���2��y��Er��3)�y�V�^Nd�X���6@ez�B�a8�3x�n��#�fMjNT�5AN��܏�Q[�[�|�SS�����.����5пa�����c֏�k��u[����p�Z�q�k�L��A�UkN��{�Ѳq��_$v_\&i�Fz=���ѯP�'�(,kQ)?����xx|�Ε �?J����4>����W���P`�&���۬FZV��HM��[��6܎LQ�7q��0Dh�@����E^�����FTt�(I�1fv-��lkmr6��F�T�8�rb�Dr&���X���K���l=����dR���T�H!�i�Ǧ�lpV�5�[�� ��h8��$c�7w(ˮ��V>q�\f
��2��O�!#�e&��=n]-��8�Ć� ��W��������{�~�^sI{ԕQK9wx���=N���MѬG;�rꉵ���[Dk�v�,M�ym&ֆ-�zp��`[$�ZV0�ѯ"��s�:%�
�=�+ey��w�e�j�Zr���/f�<��WuL���0E�a�/ͣ�_���[6����V��������r�t��\$^�qƤ��u��� ���7v�#�Z�ᣓ��<��i����iZ�a���I�t�H��o�������$��~�h��+*� �a_�:��d�]�>,#���ol��`XW;���)&�cE�_L��gD�z4b�K�����HV��a�Prs�۾�q���"�ɾF�j�C��VTG���_���l뒿��a�O`q`��0w����ъȬ�#mU0�9�ǀd!�s���Gx��n�H�|�,y�a��<O0��۰�+�P�^�Q?�D�g�ܵ-ĒQ�<�s�q���W���(�o����8�x�u�ZOo�?t��f���qG������,Jt7��i�Ʈ����$��E���'�T��G�ӝ]��B�"����|+�z5�2)an��Q�U�5*9��t��ºy=�n�3��d3�%���O˖�orW��j�z���Ĉ�"t��%��_����Y��zI�����m����_��)T���!�YL>�o�
�΄7	��ڃ�Kl�),�+��c��R�ud�E�&zX�3�RK��)��������܄diY��_�
�PM����1���G�*�����!�h����(��fOJX�������+�W'���|��ws4�"�;y&�ow驁�@x��f�y����	p�g}F���_��JÁ݇��PL��jæf%R��~�;[[;(	�o�"�7G�;�j����:/�>�&
��i�Ŝ�H�W�[F�Ѣ��mW������Ì��\J�)��"�-�+�I�|T	��)�	�o��8�R�G���6���Ԭ�6H��a�[wSi���e��)�=�h�L�w�`l.���β 	��E�s��'Q���G`ވu�89��)��6��l��$=��4&�v��8Af��2(����O���
v7��λ�����|pK�S�hB
��Z��H��񶲑D�_�%���6(J�[!Q!O#�-	��.�#��9<����7��b����y^������{�0}�"}n���`�;=�/�bK�;~��\�A�#��"�i��A��/6�����I*G��
V��e�GH{z��²d`8�z&٤��	��C/}��i�а�l8ח�WBD/gCny�o$MwU��+�
�j�'t����1�����0���%���$1�J�ʘ~ g�W�_R\]�)i�]��)�
^UY4�6/N�w���8��R��R�V`�>*+P��HЕb}������p��Ճ����+�� ���@�"��q���̌s�>tS�F�a�h���}�53D-v�w�/U:p����ҬUVS䧠�]s���'��2����['Z�DZ鍁�.�2_��VPU����8����vp�(��;���������!��bL�t���ͮ�a�x�����d�{F[�:+}��񅏟��*.�����:��H�a��W�����^ß���+���>%��h��K	�l'�Y?���Y���i�gPq�[�mRn��ݒ@v
�'��ƌ�����֨D���L�I�Cl�PQr��9~̺ �Jj�[�e��&��,SJ�.0�9�����.��Q4jX�S�6�lX`������E.�v��Mq��ȔKͥC������*&e	Te��� !������?[@�M��̿lk|�'!<���`�4��
�*j6)p�XF�/�I�����˧��R�"Lq��K/o���
�U,��<�+�$
U�)sl���D���Hf������u�'l��ӕ7���z�	��.喂���H�X�x'���H��u/ �l9ـ�.�a���T�* h��'\�8�3S%&_0B���((�.Jz!%�ǿ�1��+1d{Y����]�©A�<�FR�S�y����0#o��H��84P�ϛ�GK�"�"c����jq�ح��^)�>���`�n"�Ĵ������3���}Uѻd[�k3��W�A=���4���Ut�����65�[�߽�������D�C�b֨�΃p1��S�б�l�g��ޞ����9�O�#��'��C����T�.ɬM�8�F���'���g
��:XT����a���dL���'��e���L��ז,�~���J%��=?QƱFJ���"j��o �m�:&�� 	�AՂ,~{O�n��<gStϔ�&@=d�lf�y���M�Z�2B�Ϩ]��KZ�J[e�4�:�r�>T�	l9�L��C��Ҧ��j�v	f�\q/d������� ql�~���Y$s6x)��7eP�d��r!���Cg�֠�]��V�.�07����0n��]y��� ܯu�a��/b6_�x{�ӽ�R������hyg.�q�jV�Pݏ��	��ʐٞ��O{�R��<��ˋ��.�[�����Ъ4 z��kQ.s{�:S��̯*T�i��`P��tz	�@��ξ��(��J����2R~�f���@5cK��r:,2��ꡓ�H�L�",dal�|�{���9p.�$m
 V#�%���.��Ϛ?�z�'X�r��[n3�l��f%\���^�v�m�2�e75$ù�/M��:�V���2�Լ�"B$����bLhY�}��k��x	�	n
*�xL��1�g�q��0��B��k��|��'��b��F�E`��z�l�I�6��ޔlF�m&z��� oۍ�k�� ���D��nD����2e��e���ۥ/ ��>�P����;�"�xD)L�5rU�.��	 �l�k�� }�l���Px���
;��h�u Y���	N�0dVv��AB���}Ц�PC��ȃ���@ԆR ��`~�N�ރ�H��t�&(�T�J⁯�Pee�u~�=��������~��->�4���0Vq�؆z�+RCTL�Xh�NL"u��S�J"�ǆ8F��U���%#)��Z�*����Oy�v���Ŋ���o�͙�����J���ص��I�C�ѣP�؈�����I�ܴ{q|�4Y�'"�Y7����o#	�&t��V�\�A�X|\�.���I�������neL1���fm�7r����B���j�\��<j\78)7�L�z��������_�.`6���2�v���r��%[æ��w�Ztm~�Oػ�Yf|��?���֩�e3>�������"#��d��Ч�{9 �åY9�Jk	R��&�d`o����6�n;�+9B/[gPy������+� �=�'Ϳ�$o��fRr�E��7;��V��`��-J��B�#��ho�,С̼��$M%Iw�s�ؤY�_9	w)��3��D���n3����%*�Mk�s>�Zd--�9lVI��.5�&r�4�[ˇμ�]��%�ϴ]=[�D��U.�=G<���:�H��B��
Ļ���#�����q���/��A`�k���Y	*���ԙ6$���,m�į e��|�?�|N��we�HL�A���yd���/����Ы<J�5��J`{�W��e�������x���~N.���8I`9��j	�Z\�׺�&�d�C��62HĪ�R%�x�K�g\��Z��f�ޛƔ�@kU�`�ǘ����̛�<��1� �@h�d��ex�1,j�$�_���)		\�c�`��N6���'���'��sa�����@��1O_��i��nf���k����邘�um_T��|:o!T��t�0U�FL0��[�H�PDK�6��&l���Ȗ��tu=]��?c�A:Y+6?�6��I�-�!D����S���L��A�Q��K��S����a?�)�������,l�	�K`dD�y�{�j�����ږ��M� ���v��.�@��������$`U��V�^��L�J��"�%�P�-�Y2cr��x��,�츂^^�5��(7��5鏦̘�1���}��?L_{|���
!��'3�N ���B^(]0-CDAm��h���S�w�4���s:(0}�0�cK.�4TE~*��e��b7���0�VvɈv[T�����:�$�k ����Ŏ�c�?g�v��gpxߠ�Gtm��b[�69���|�`���Qa����Іt@��$[�j��y�VZr7�cM�����fUE �[��&0�dwd
Y�Ƅ�LN� \����\ˍ�+����"n��yTE��R�~�[#��}�m�"�/5����_._H�<{f��O}V�y-m+3k���B$�����o�0�J#3inn�G�F
.���Btӆi���	�q����<<��`��e~W:It�v(��]�1��8<�)����D�"���l�<�.���P=��g+�m��_a��FY����`}�B\�T@.�nKʢd�\�B4r��!,(yր��g�=�h#�$H7F�#c�n���fK�!�(��n	�e�?-��2�;n��ef�ߌa�T3K2}������
�u���G��b�f�΁�e�"J?���%"�V:���yW���Lr�F;]�8a�����x��AQL��X�Ψ��S�DK����
���}�4	��^�:��=��ag��uo��+�.�� ����Υ\k�cY���wj=�N���Ũs���W���je8	�l?�
�}*�2���I�{�����#�
�%%��T�5s(5)�kY�����z�N[~���p� %P�C`[�iS��QE �sxj������,��J���$��t��u�&G�i��P�I�(���(d�'�����Q��TF�%�E ��B;3���<����c7��>�)@`���Q�%�:�@_� ���,�e��?�ڬ.-�ڛ^G��~s�\�]���=�S�[���dFCa�A��)�J���V�$q�E��[����X�n	������k���I+�B��D�\���k'|N� ��t,8ؓ%�
\<:�k���U�@�Yl�����Ǒ`-{jV� �{W����23{�x!A�����C��Hm�����$z����76F�-��Ӥ��е_��;�B)u����&%l�$V�X�B�����4v+�O�<���~E(�(/[�0]jAʛ�������+�����N�+�:c^�%�~48��6��,���ݟZv��s���A��~Q�a'Q-�Wj�:Z9��ry�b����f�{rCI�35�AÍ������?7W �k���nl;�=`���A�����e�4�<͛�M����@x���	��q�����W������z~���b-��8'"p��<��E/U�5�Yj��ű'�t^l��	L��C���h���v;�C!�豣@]���mħ4w�^Q3� �a��9{��7��2�'x�uo��0벯�H�O��]�Pk�\�� %6�鎚�8.��;c�0��/����z@�w��.pP�9ѧ��:G9�����+w+s�!৴��֞��:F�Y$��|��4�����o�n��K��Rewm��k�E5x�$	U2��������9�RƐ�ߜf-S+���(�@g��XW�=�e߰'*ds��њ!�� �_���o^8Tb`�B1E�?Y�j�vz��ւ.��;"�9n6���x���8b�p�՞��J��ߢǓ������qX�>��잦2xm��'���n�0N!���|����'K��_�(q+Ů�M�t������~��w|vK��%�
jU�y�5x��F�����Ip�Ei���/r�ꅚ]�Փ���%S�?�5Ce��p��}j<�ùZJa"��2�z�}E���������>�{?��3U���5��6�Ja�@������P�^�廉ͼ��P�G��zoIA,�su�N����Ʋ�m���Mu�#b��ڟzM�a挟�e
r1�K/�r���or�ާ��2����!����C�	���{!'�C]��T.��$
ۺw.l���c��Og0҅e?�xy흜�io�j��[��1���E��L�MxZ�<[�*PD�v������|1/.���(q�د�hi����ĝ�0���#٘��hν��#XY�w$�鶊���e�9�ZjOe-	�D/i1������/Ĩ�@i�	����s����7!Q�߽V?��P�<t�)Ӱ������g��4���!34>V�G��d:FZys��ćNBU}�HĈrq;hªAH1d9llr������|���A���F]��T�WS]�I$춷� ��&mO:i��N���U�`���� ��Mюe ����Z2y���w����?II4н���7�|,�.}�:K�*�����;��J�WK���\.���W�x���#K4jCbSyt�̾�'{Ÿ�[���<�����W�.�6%9.a�?����6���`�Vg$��?|ڕ��%[�i��?A��L���ϵYI�Pekq���]�2�/#���mn^��;���r��pp�������»=��}qB�y3`���F�Ġr��w�)>*�acp��}$s��Wɿ��ݏZnfpbڒEF�ˣMBm�`ڨ�ܾ²�{�q���x��!"�o;�|�s�Yv�����W�q+N���B�3�x��?��������J�ve�j�/B��J�_�Vܾ��Q�Z��Ϳ�*�7�xO��x�C��ꆕ �~��jh)����d �
�iו�^���-X20���L�)vY�ֳQp��J����) ��$X�Y�Zԭ���pA��	v���Ti ��a��j� 2���L�f�f0h�zb.oT�֣�!�Bи��yZˋ2o�#g�ڣ%M_A����F��ݪ��g�{1�����j�,Uxy}H�x���z���Ϯ�3�,l�y������EԸ�݅+Z8FuO�ְ�D#�:�ti�#�;]����@wa���_.�7��GZ���`]cA���ѹ��tF�7R��f.�^tɒn��n^�!���طb��)�&1!-���}�廋'1�E���E&��Y~�j�،�p���v	4���<��0'(�zç��0F
q�H�J�g����]�6��܂��/���|��2z��-�=���/���F#��B�F���,	}wc.2��ׂCi}�����'��1�����p�'�2��<>��p��� �{�3K��
ђG�3�}U������fх�K�Nz)�&4/=XԞ�d���7�»z�d��oW��K�s�	.H�XR ��������,<g$*��U��Cf�Ke���n��}9υ_R�z�d�&�P���н�q�d5�B����æd��t�
H4��7��Y��6�e�!S(ޚ
����u[�`[����{��?5E��>Y\-\�`l�'[�H�U���)�t�������]�����%�Hw��=���y$VՏ�2^M�GjWL����-f�܄��� 3|ة�����ۿ:��?���0P���F^{\�����s�@����mb�d�ڥw[\��9g�)v���c�O�����F�>�cͬ�����:H�f8wҮ������pj���G���tO�R�Ң�]�<��w�I��ˡ�ٱ��'<1xU|�kd2иY�z�B����$���3�׉&��i`,7��L���Ùgp���>i�&{x��Dނ���<�8)yM�L*�uW�P���9�������F�|���m�x�<��i�+x�7>���wD��/^����x�+q�3�`�˨ojJ�_Z��pV�D	�X���"��զ�'��u0.Ѩ,7�Bf��%x�����
��W�O��M-��׿�!��E�1	��Gj��lHd�O!����+��"��XG��徴)���`t�*��F���\!A���c�}�4VҪbt��m��y�Z��	-uS���I�OfIcS1�w������"�4�r�#ٲ�Q-T�.q���푏l	O�S+��G��h�5�7U�5^X4�K�o���JIG	�;5������#�����U�
���0!�����0[$$�|�M�?��m@W�g@WǪK,��0R)P�F���)��?�VH�o����6��:͑:T;!������8"��
�,�1[��*���Z�4��)�AK8Nf_#���)n�v��ξ������U���*�{Lu2b���L��8����By,�}(�*����m��4A1@!��3~ɑ �s�@[��}�mr�X0Ww2��dz��+N������Vmr/h��LY�l�%`�CiE�F��2]������!��7q����_��N�����������*���j���O�^�����Y{�͗�LF�a�]��[����Ѹ��ϦG�����4�Ĉ  s�d(�A���/(���s�q;z���y���A&8��$�a+����l��ؤ��ϵ�Z
@�����Q4�����$@"�$5C\��՞q�.�M�ݔ��$��,����M����a�/dmx.=���-�ow+��K=����o&,C9+%'4�E��n��yAZqxm�?�h0X�7�ݚ4�،���d�D��W�ˠah*�Ȗ!���	D<����(!��zB�����y�)�6k��(]"��@�Y�7Q89��s�V/᭦+7��#��6�{���%^y7�CZ�k�wT�����
������xx��g2��;�`w6-�"�S�e�g*����xe����R�}*��8����!��p	3[�y�.(��d���{{�*��<�t�B5�P3�ٯ�5�,V
�� :n�x���?Z��Hp���+���ߡ�i�'�+v{YA{S�*GƊ\���Bj��Cu5흝���?��fDǌs� ��8�~q�/������� @}M�q7��|�oe�'ؐAC���l�I+�#�#�I�}�)�) jG~�4��u~�8�O���)�Q�#����͚�&��0�;D��>�ٮ���#�`��3��� ��1�۝j!/&�ΌH�8��
1ԭH�$t���k�'��.(��:�1;K�Z�_)IBx ?��}3�/��ܔ؋�/gR<��{�#���a�u��Pc�<x�n����o(������V���_�/����^\���Y��ܶm��G����B&3$'M o6�<�.�|9�w�k?֙���ug< |y��Ղ���iZ�Q�c�61 �Q]���Ry�ZRi�'XB��,�Z^�;U�Jy<�l{��	{�f���J�Q�*��E��5˓�my�{R���NU���h�F}�#��b�vA�*-`��t��/��h�/� ^zZst��k{��v��h7�4tR�D��s��_��
.]��� -�q�O$���f���`$L����~KQi1Q�]�}<
�*�����
4�귚�Ⱦh��-B�����=�_W��t�)��^5�]�#�y*Ↄ��R�9mtt薉�{�Kv_�d����T��P�d�'�`6�	�1V0�\���q��quP�E�BwbZ��l�jdчn;���[��1���%����6��t��g_6��&2�"E�l `<*ů7�
Rnn�+S
pKd����J� ��y^D�	]/c/j�C�����@���ĳ�)`W[(xQ���u�
��Mmq��l$u�^P���YR�G^/�R�B�#k︟���V}E7;�nt���eG�����5nwd�H¹l?�Y�j��إbS�� �h�O
�.�tw�nwÉ��r�V/�3�ˌ��9ѸT���K|6��ֱ�zgp|h��"A��n`�LQ�L|�_P�Fun�E�Z>��Ww��AȝN����k�)�v���������~����Wؐ��Z�rT�=]ܗS�RN�}��+�Y�3��`G��:�?"��"�M����c��>��O61
_|H��PZ��ے�g\�4�������~���^R�W�M�xAj/<O�a�|MMr��h�����Űw怩5�7�7{i��R��/y ���P�xU�
�4��)�+�e)(�	Љ�*�ڼ���
A�o[�0����$��Q�ş��Y��*iɚvP<��YC��	�ʆa�ս�7�/j���^T����,���-�ː0�8��՛	����B�-��v:�G3k��V�%gk[?�h
J7-��4�ļIu=y��y�[:��x�o�6~F�박��!��;)��^j!�=ѵht{ ?�����8��:+XN�9�1%z���,3�?�+�G��Ȱ���Ħy��*��w���0��
<�\ ���A*�"�-��Z����5�51p玜��Q(Ml�|��D��SЕ����8�(�DuC�`�� �^�^�b�$�/c���!��⛠6)�uU`JRk���H��d��~�WȖ}����1 �˽V|f�}�ⱴ�����>kR���*��\�,0��v���@Bh�O6(��[rz�AILDiG����\�h�(OH�k�C��E�J�B�(=z��w�*�O��[vRʬ&�k*� 1.p�X$V�])ؿ[L��ߗ��� �]s��{F������F���:����NHg=�^	�|$���$�Z�	~��@�\�/��|��G�P�;�Ǌ�06w�����3�7�D�7��	9�R��vm\*��_mz��T��b�M~ܪ�pL�TĶ�Kc��vׯ�jc�1ܼcW��M��û�!j,+ w�=~9K(����N��4��feu�ODE���g�"aOgLs+�ɯlt�H���12��?��R`��Ϡ+���#��&�L�]K�͒g���\��!>�@���i�����e� D>$s�2z�ť�7�2�2����^\he2굝�>)l��ή��,X!_�
��H�Gv�Q�ηF�r���v��b,�#����3��}���Q�ҬC[��B��Up�x�\�/�3o�$_hK%�����L�_	�m���l��"������7�Γ�JL��.�?���n�?� @�H	���$>i͇�TУ70*���?�j/'WtldP��#-7��*�����W�6L�VOU����P"��7����A��h�?��/��A���%��4���>ʬ|Gk���s�ר�����Na��\e��st���%�Li&�5x�קk(�A�s�^`g�*[n�.�V �̑��#��7)p��q��g�hP��)j�Y4�N	�[+x��8��LPB7q�T�gEgF-�u����y�ȶ�0�S'6����iv��
s�����G��JUS���-��È'^��m,\�S�\�| �*]�NQ]��k>0a>� x�d&��Yd����!Sb�U=��"������m8���#��Y&��H�
�{�n�}�%ޞ
ʐ��h:�.yC<�w-�k�٘�_��&f��Ԡ�Q(���z}��?��Y^��#�q�ş�mT<z��3/��j_��`Y_���С�I���G���8��2���Þ��ª��Zt���7R0��"��ݎ��C"��U�%��y����O��0��g�Q�P|/T��r�rɔZ>�U=C�~)��I9��\/��H �`���1�~B��h�k$����M�V�BRR	��|�5��]KD��!�0��,�&���H�IVڦN+OS�'H
ڙ�w����2#j �j��}�|G�����|
ҧu]9��J�x��N+Z����
H !:̵�;��/��I�wVh�{�e�����Z���G����Z���+��M�."4@Y�;��?*򺎟`���9,j��|����S�\�i@��w<��=�9#�9�+4���\�df=_�� ��n��8h���]�@�u)z�jT�u�/)K���u��?;�pZ�/���^����q��S�V���E��5�_9؃���"ā7 ��ـ^>��G�)PW/�0���7�륄�CMb,�	�� T���%��/J�0�UF�
!|s�ﺎ���n��]7y�_8<GS�A��{U���sJq���&���.�(�J\62��M��'q�V���D�C�A�m��f̚x������͋���>�O����P�62�N�\�='@V�z$BrL��H�<��:Q�P�n�j����7���:�M��L�,��t`c%�sD�
5ǟ<�����H��5�|��se�-<|�mv}���6�����˒2g�W9���!ݖ0��eJ�)��Aq"�KY+,�X��"�a\��{7�D7!s�������T�/�	=�av�,�˷�m��Vp�n�e~�Bq4��I ��k.U�Z'�-�h�Q�Q0͊��m�K㕧SW��l9���J��-#�JF�x�і��~��u�Ik�HKX���7ܝ�L�q\�n��5 ZVp<:�0=!�:�ׅ���DyG�j��H&C\ǖ�̧�k��3�f�ڰ�5��7-�D�G1������Yn��Y� =|�Ü�g>w$o�4z�hȯ��J��Ei�n�`8r�����G�L�X�bN�}��R�]�<����+`&#��g�IQM�`eY�,��D��<Ȳi@f�ad�Q�����c8ڐGv�-��Y������P��|2�������$`�N���.��$��K�}C6������&�s{��
�eF�����+D�s��G	��Y�4��fH�P.��gƲ�Aj0�Y&z�ܩ�3���]l�i�Tx�]�����pќY���*�`)���ᏰF~������H������z��� �,uۑ ��B���!��O�'���3�G[�����_q0񔴻a ��'n��Š�[�'�iߖqv�ƥ�:��8z��0�|)�r������*��g�OLo��+Kr�$F�d�$-�ӓ����o�z�Q������z�	-��;�9,��W�|��̊D�g�Y%�KL<�*v�S�2\#l�n�7� �Eb��W2�~c�zOr�$ywҡ:�],�)�h��U˞�"s{�T���h�����O��Ƒ���1�x��_i"�[e�;��͉�8�a}Ar��whu��\�&}�e�T��D	؇�1�o��l�v�Tg�@e@���<7̉/��@RT	�믱N���T�J
�������2��_E���U��9���fk�W(���m�U��������ؤ5�0Rz�ޞ�α���ؔ/���z�o����unuK�Ww����6��_�P���5��]�3�LLU�iܬ��zcN�u���5��:2�LhZI���4�L�w�+A_�e�#�j�E�����;�?E_��ʻ�Wr8�>�$xu��٧H�x�,�U�9�j��萆�Wt4l��1���ȶ�I d�	�>zW���5hf 9�=�a��w�x%ba�;T�D�,gT�f(�74�aaL�M�	�zd���rPSm �X9l%LO�쮢� �Ce��Ύ�
���+(~��,_�I�S�i���{*�d�|����g��v�]��D7�N�Ѣ�����QÌO%h �7�5Pё�R�pp�b���Ɔ58�� -���`�i��V��7Y���_�&}��N�CU*�rfL�����3�V��]+���c�kcc���;�{�ߌ<����W�
�c�H1��j��N/͌��8$�]��@�%Dn������x�5k%�g�O��	\�z�lT�]_��W��bq��Էd��?�jE��"�N!&!&e���[�j<G .�뉩6��E`F��P�!SG'��TR�X��7���a�c�9�����#�z�b$+�~30�w�,�Xؼ��2*ф��\	[; z��s���� }ن�5��P �2���#�N�حQ�_2 ���K̺��ɳ��	�N�u���1���j��R�<6�*ؓuC),"R*�e�ί�̙�y���y�������;�]������|Qu#������Q�v�"�_�t+�pF5"�C��mg�_��_5�Ko��˃"'?<m��<ޯ��L��]�B��gf��%��m ��8��и��6��D)�����r#�0h�\gY�����c���[M�?5���9ޭ�TE$��㍫ �\����F6.e��҅e���9zl��m�Qn\і^ɟ�Dܸ��b9�j���<����]�߃�g�L�9"��vI�#��қ`������^	}w(�`�Z���c�����	�������=��(��b",:Ӛ&�I�8�/�&$�f�^�A����)��5���[Q�ލY�@E�̉��E[J��O.Iu.��z��Iԏx���,����>�z���d��6x%���;��������DI��la�FD�o	�~�£9-0�W���b��f���ɨ�u\/tu���.�.��(TTv�\oA����؁^#�7�*Z�S��C�?��)vG�:���WЬf%ޭU0�M2������*;�.g��q�������me���%<b��)�a�xʹt����Y@��$��X��0�Y&׿�1����L����@q�=͕�l}��*~Ѐf��4�8+��88C<R��w�a�L�:��Y9!n
��٦����F=*&��ؙ5���ǜ/������R�-�v\֟ ���hl5,!|xg!�@z���\�W`��F��Ay2�Ώ��~d�1�[=χ������3Eͳ�#�qF\�?��k����Y.ȋ�|�5���:���`q�W��t^^�|�wR����c#?���Ba��K0!�T��G��%#BC�u�W�s?�����B�`y��9�CX��W'���W�IԒ�}z^��s]t�2S�,_��2�Kb�^ά�:����F�Q��
�oX~
��Tމ�K)�%���8�R��'i�4،��l��7�8�Pܧ�Jp?���E��Y$��	�D��u�U ��ɪ���ߣL_n�m^�s�OB����6�Fbv]I�0��U8�桁y��Y�OУD�RN�N�b�+��͍K��!�|�<Y��BR�C��r��b�+|(������t)�8�Y}bj/"�	u���`��Y1<D��y��(O�7��?'�?�F�8�	Ɲ6�Ң�����f�� k-T�]�w�_�]�Nu���NX�bቤ����4����G�ʆ7!"M�`��8Ԃ�n�6a\+�vġT��4&R�H�~�

�x��L�N_�:���<y|3TA�霊)�^9u���d��+�q�?O򴍧��}?�7V�к�7���z���tP&��s�I��Td-f�xby�m#u�F$F����;j��l��2�ⰶtq��2��tJ�(�Up*LǱ�#761��W�}�����Y��:�U7~�\I~?+K*�s��͋.4=�`!�j�Aj���b��������N�"�s�QU�j���������b:��D������쳅T���N5 ]��_4��%ߕ�x]�`n ����I�H�Λ��|��j�,�G��3h��Y�5HE_��൴�wQ�pr�� C-��׏D]r�	�ſ;�m���o�;��a��~D�jY|��=hm�u�y�Ӛx�	�X|\m����+�ƤB˟�� i�ly�c���Xiǌ	(@4y@��)�%-�XWR4ݲE��\�¡������-��1���/�)��%>�ʟ�g��=q��U���&��ggh�l��I�Gn7�c��l�7֑7�k��j���2l"�1��Y8utosb���O,ZaS�RL��"_��S�$O�)ї�z��z��o�n�^%}f��6AOTC��+O14]���*9Uv�a����6����/����Nԧs�"�����¦�-[x���{3.E�C�����rFX�S�%�����y~�{�'Ͱ�#�[T/�d���|(������f:/���M�U�?o���+���ŀ>�H��Bx��,�cđ�(�:�v�>[iH.�Zþ�D�*�i�q@�}@{�ɧ���Vp_��V@C��d"D\�����J��C�N�c4��<�����ɨf^<�$R}e��ͽv�%��y��\���F'� &m����3���es��Ab�n��:	�,ZGyb���W~�v}Y h,��	?����25�����v�K.7��TҦzܮ-�����A���R�%.��C�������^��#ϑ��.%k<H�vxL�bVO�7�b�?��z�u��9�w�Fr��m�P�z��c8�*�!��l������MO��N�F�C�AT�{F�Vf[�k��a���;��o�fjRw������v�1C~�)ty��%
~T��b��Ί��kz�s���Mvq�>� �i�cFxe��Y�r�4��j'��67oop���'�7��kD��m۪H�������,��g�Hm����l�V�m�{ܘ����bQ`/�\w�ц�/�n�gr�U{H��R2X�<w���A��d�>�\��$풄��,F���E�j$��ؿ�)=�\����v-exAMV�+[[4D���o�(ĸ^�E�5�4�����v�ןz�Y��÷`7]�k#a�(������W?��~�c������r���T���d�-	�ȕ+hOu��S�T��a������h���[�k�E�l���K�v9#�A�9�cJ�,�s2t�o�`�q*��v����3C�u��kqZYEƊ!�������?FD�6���84�5$+9ϓ�W-����d�mZ�GA�p9���=��w3)��Z�
�q�Z7?鐂��߯;c."�0���#�#�n���<i����nI���"��E��f�ҝptó(���u�iz_�8������������okR@�!��c�^�b�Ͽ}�]�s[�}�ƪҲ/e�p�p��ķ��o )08�]M��0Å��n�\�M��{�,H���p�x����#C�B�4,�.�u�i����1/��ĿiC*��"�Aa$�f>-^���"
��X�L�v��2��a$�y*oV� G?G�û��k�r<��'�k���6Ǌ��R�K� O�[r<][�t�M��V���p����F��U�0��=uRV��6z߻@��u�^�)�
kn�vq����O���O���yvK����,�wH��t��o�^J�~�8��\s�IC`e�š�_A����x)��+�x���f(�Rڇ-Ǉ.��qRX��zQ;��d�5�|����ܐ��@���Ե��o��G��g�nCI�6�JVލ�n��ݦ��
�^�-�hH��N,e�Be�oY<��zb�MWL�cN�uܯ�7oAK* ��2H��P����L��6�8:���Z��>ۂ((�&,�zP�
/�h�:�8)[��DR�)����ALAa�CВV��!��\�������-���qB�m{����1Yd]g��*M\=��7�����O�"�DZ1����!���_ѵ(dT����!�̑����S��R=����ť�ԛY�Ҥ� &r_�P.��dĝ1�"�����e�&b� �*ys�V�?�ό�?�΋�%{�_�1HF�h]�ak��j������-W�˫Y2��Q�ׅcI����8�p 7���4��^�b�:"p%����sx�o���9��Nj|����*:�c�7`J��c�8�|����8V��|5���w�n�H?i4T���Q0��0���O���I&�P���Q N������Ŀ�2���4�h��h���YХ��5�E�3��,̦&��-V<����/��Nrɡ$�^s���^���*���zݓ��`��iZ������!�ڼ�Xb�����{�E�ѣ0�
t��,��؅�~][�=_�W��DN:�V�}F�T��m�@��dƠG
���������x���z�X�t��R$��0n�A�`�IZPaI�ᥒ	�9.��gW=,<�R��ڳtgEx Y�[�����I�����4WdL���<$9���|�W�7��	�g��k�'~3B��ʮ�RQ÷�3#�������r����<��N�!��ة���;�38@��p�w���z#q�����{�< (S�tr��D�� G�!@΍�hf��V�b��@5�[���($������[�S�E[�Cy���ڒ��܍Ϳ}`�Q�yf,a����Rz�̅�j�]��;"n(Q8Ǩ�Bާ��ÍRFяaM�5��i�?�?#4o��W�F�㕼B�I�oa�����$M�AN�IA(�9�]v��q󼯆�1�$?E[i#:�$�x�������Q���+^�x���f?ڨ�OL d�ZG�� 	<B�ꭇYL���г��K��!O2�E��5kX�c��}X w�|�+@]}�����p������I8:�D�ux�0�%��8��b��șQ �#�9cҽ���U��l�{h6Ei�	�\t�R�5��7�̗1ck�z�Å�e��ȼ���<OGY���P�� ���Ul��7$W4�34m�$G�V*y7�:�"x����י�Z瓥��[n|���y+��Rs��O�IĻR��t�dH�[l*^m�O�Kԑ�(N��Y0��-:�v�,i�N�(���.-v�R�M�t�p�̊�T3�뚀���=��}x`Y�j���b9+�����F�c�F���%s
KyE�!/���tj��Ö�Fs��D�f�Xz��ӽI�V� �*?�U\�e���]�B��m�\КݠH�L��:�o�P��>tU	Ϥ�ʎ ��䑏	Uǈ� �����'5�D�U��;��Ȱ�/[�U�� {�}�^�Z�`�m�t]�w��E$\�y��ί�e:2���ϑ1#S��ކ;T�x=���#UM��EC�r<�ְ����T\�����S�FZ�q��	Pi��G�/�Lj�τf���t� >�"��xtH(��r��3*��n}����r�|��� &;�u����r<�o��"O�x��T��!JgSWT�sZ���`��Gα�ڨn�[�9H�P)�X��%R��k��O�MÁ��;����6�iS�9(k�\`W�[=��Z:h�<T͗[^v��~n<�b�+yDú_86�RS1�����&B��Yh��B�
}�`�uoeH��8+��c]�/�	$)����o�[۷��9*�E9�5h��5��g�],\T9�^�l.��_3��-���)[�wq����p[U?E�R����
~��S�\�w*1�q+��rd�Y !�ėF��`%~&M��������F��%/�4tE��f�.��X7�3��1�i���I�?0LtB�m[/�4n�,L�A9�� �_��!<�Vb^�3L�B�f��řJ�;�t�KJ�h8�@�{���3��"Hpf�?��wb��t�ރ�'�SP�EWR�l�Q�i�'�("�R�~!~���E[�{ʻ$�SO�����j�9?�u��?L�Ved�u�\\4�':��xA����PYθ�a�Tz��g��̅��8`K���
���*��;^}]��-b}Q���*!s�Lxҥ=�_��t_����/Ǻ�?�bN`I�%y/s�-�	V��-�~��������Fׁ��&�����ꢂN�z�_Zv�buU��bRm1� �]��$wwwL������z"�>9�V9T�i���b�4Ԧ�iR�xĽh����>e��%g�"�	4�4����������#���X-�[�(p���P唠@����ݥ/gm��$���z��Oe!钿���%}��ҢV������>��ꞻ`�~���1����k��~�r@�d�(�Tu�Pe�p�&>3V�؀i� \H�"�t\�KE��Y�;\j�GQx2��MNG��1�	X������h����^�mt��h��%0���r�R���:3+���<ި��lK�c�	1�x3<l��s%�#�ޑ�U�6':��2��u���N  �&	��[�ϴ?U�0��2���VjQ�)_��z���!{N 4����$����7�� :g���~�j����[L1�:�Zj��wU�/jJ��B��ޝ����^ܒ�:���PW�o2���e�ϧ$!ZG�˥F�h;��%滴�k,�07Ƴy��;�e[��ֶ(����P1��UIi�����0�/1Whb�$wi�<Mc��q6�9^����>!n땍흥Vt`����3e�NK��4��ЦK��������+A����`��X��#,�{	U�O�OB���f���!����x,��d�\�/���S�=T=ǝ�Qx_�a��$�5-1ӟ:�V��Y�Ｉ6x�
�Yq�A�ZM�0��֣���v��e��Q��T^.6��P� "��e����{-��^.:��D����Nśu4�Z��f.Y� ��.٥�D�D��:��@��.�V�{�P��,1]��r;��/�d���7re���=�9��"�N0�����[���M�/[:�%q�w��e =���Ծ��3�5q��:`o�<ߥÑK/3�	2��n���"��)�0&Y:�?L�m�XϤ��a�&d�Hq�~��)��]�R���i��=.��K��x�SV�Y~3�6C�e���ȼ�̅jݣ?��m�\��G�� ���h���h���TE�!E��R~�ߋ90i�m.9�tI8h_l�6q��D* ��bH�����@Wb�
�eR���[���V|/~/8�BM�8�������פ���L��y���,��2�����Ѣ�vn\��<BE`;P��^��_=��3�_g�)��nY
E�Dc?T2�?�����@�ٷҸ}�EY=L�H�F��pg�͍���D�6�;�b��om��PT/�H��`�,�lه�!!��,�i��� *�pХ�,�,"���)�����N��B�?�@�M7����K�͞��I���"تv�"��C��5�)u?P�HA$"H��jt �z�f�:�m������C���<���1�ȺaJ9yq��P���1��^��b��tn���u,t�w;/b��4�2dH�D��6�6�Ʒ,ٙ�r|sKQ���3,~Cu��z��A�[������!�ԫ��i��E�Y����y����+����"R`Z���tִ��UÞG���;$N�ݤ�5��%P �ݡ������w'@f��!�!�''�~�2"�kc>��,&P��3�0������W��y&�Y�k��a ��v�H^�]�sɧ������T�� ��z�?�Z|�y
�rT3�1

ࡅ�&g�;o"�"b����1p?I�_�w�SR���碧�
���z���D������rm��y��zIFP]�` p�Vy�TF��):��?�����! ;�g�Z�F'jKۃ{��b0�������+���"+AYo10^�H��DK��c���.:%���rh�B�Sz>�'@o&0X�_%F�8Nt�Qc�Lh�h��󞓐����J�Ѷ1�f����jQX��!��ު�4�������!�w	���A^rG�~Ӈ�z�/8
�g�
�;�.�K�$��o�( ;a��LkyVƑNI�vyֆO�ML�:�.��}-�iR�II�v�U�L�)�ޥ_�%�B~�bP �dDauL �#2_�=��?��=��`,(r�ei�Q���*�!9���m)�J�䂙n�)8�56��H��On�~�<���5�i�:��ƻ�z���Q���n ~B�\ʌ&���jyMJ}O\+α��-t�nܖV'��T����Z�g����� ��c�����)`�+�m�z�ݫ���6� �1����W�����g��B�jnl�����A3��AK���$y�v�k�]%��Ay	l=�KBo[c�@�FA��a��j���('�P��	/�(
�*���,��i�JVe~������L�ol����1zd4�p�Z�jP��])5�+Cݻ� �s��6��{.�,��%�-�+)��d�\���@+1�*t"�����u]�g�J�M�C���+����P� m�}q�]ׇ諲������y�»��(�Pd�b�;*���F��L�-�n@~9�*� �� $1RpK�������w����~��Lz9@G����� C4�v��"M8M�']ro��q<Ş��i�5"Jz��"��Ac �H����d����l��i(%�6��r�A2� �9����q��1�T���iR�s	�i���G���K�=�L��MZՄ�Ve�+X�?�3��Z�;UD��i��*�	���/L�lh�Hˋ���HK9t.d��� GEmy����9�z�3��;�����%�_�;���+���`y�=�[��m��޿&cR��0K���Ru�v��x{~��;ډ3����r�! �\�jm�����*���S����jI-N�\�C���i侒}����n�l���DB]���'�WO�X�1�l.R�$�.��j����4�		����q������t-�f��������J�V�{��vu~�������"��~���F�>d�C�������=NP�ZY���Y9`UR��y��H���Qy0��@�AB����+�������`��r@���ۭD�/�۽\�,)K��5��h�_hw��^S@��c&�&jE�Dh�:�'u�&�����U��ÉY�@��iP�N��ǑG$+ؚ�յ���3u^"�av8�re ��!�1�/�6\l�<��'�;˚Q1[��Ӵ�b�]��~� ��w\ɔIw�VK����u�������i.�Ի���9�����@�{p_ٝAF$Y��z܀��6�!�N:�j��<�ʙ�y(	e�K���K΂�E��^�ϱK+����)sq���#
�M�VPK�T��YB��g��E$�u7��_nrmq��̀yv�P���wV�;3Ѐ=�P�w׍�$#�5��-ƅִ�S��������	��>02�c��dw7`�V3���[��",�8V�k�R��F�FNf o���2.�b�!��1�N�=N^��H@���.��Q���D`�ܑ+�9ZL6�b&&�}�*�_}R�]=Y�!t�.��jKd7�e�ՋӔ�nLy
:h��sHҵ���
��	��mNwN��O��b��Ǔ\ Q�96��pЉ-��ʍӐR������goM�Ioڤ>��=@�s��1�����ف�(e��.|����,���늎4%!�Th��ս�w*���Z��ɛx���3A�C�+�W�b��Λp�
n��^�e��g72݃�\47߰6%Y��o5����s���'�Rd���4�B�%�o�.@�/���y�����
@!<����|~Q��K�����ţ"���� ��)�^"rՔ�u0'�b�,�cEWlUcN����#u(�[m���+����>ߙ�,h����vU��.*�Y��%VR�s��G�B$�b�B�+F�	f��Y�L~�U�MP���A�w���H���7�����M U�.g����1���((}3zѯߴ�)�j��-��-���fp/d#�.��I�m��^�0P2�_]�%����u��z�=(� %�5PS�!0g�w�E�<L/j��2_�7�	��ED��ڠs�uV�oqt5R$cm7�UOor�}{����M�@_x��D1o���x������(�Դ�ZO�tI�q����}�,h�E�?�V���4!�d�駈�p�,��ֳ��F��k�u�N���Q�A���D���I���{�V�4$�B��� ����7k$A�xFkv�ņ4 ��N6� �}�ԙ���9�+�C��s\�����M��{�B|/*��vO2�ڪ������ǥ�1���3���<h)Ћ�(&�?#q��U��M~������7���G5�DS:u` )�ej`>	7�i��\x1�|�n9��ź'�,��n�G��)�F��N����2��uR�f�ٿj��c��\�Ag�3��[+`�9	�$Fce~8c�H����Я����{R4N�f|r'�Y�|֊~q*�#>�q��M�r��b���4��
�&L��Q�fלW^�T��� p��� ^O.q�������H�~-��ᆽ�3��x��j�^7x*F�+�7�2A�ty��ĕ�E,���6"UO9-s�e���y��چ�P��%V)�ao�ԋWs8_���o�z�z0���OS��c�w�D�o۰"���Ƴ|��-*�ށ��ۻm+ 6���'�[��1)w,�+�*o��f��t�q�L.�BE ���يP�_;,�{+O�$`<SD:������'79�:*:P4�BsDbue�9�)�E�`sѭ�^���Cb�k������7^�j�t�:���}
���~��:ޙo�dŰx�P�8��3!J,۪]�Q�hɷ�k'�]��wCs]�pڢe�A�E�2g�d\)UkΧ.{~��"��~��ߓ4�M>x���u��.RP��M!�j1�Jd�;��	s��\�����4M�����)-�ҵz�\���j�߸	V�¤��Q˲���]��6��tFfr\����8��e�C
֧��|��m�q��I���vԕ4�EE�6��s/>�q�	��l�z�m���.�8�	xgA��	ޜo�vv�rd��2��T&��Mz6:��A�߹rwܓ��&Ta��mV���
���p$#%�y=6#��)��*�yhKp���=�ܻU}Y���CВO��d#QyWI
�{�[9 �T����=��V�֜j}���ն�ei�qV/�L}<��R/8�q'v���?�m�3ld'
�ԝd,j�.7촰j뿮�W-�0P�H"�"/t�j�{Ґ�OF�Q[E	+�DȦ��V�����Xό����+Ž�q���~�ZO���"dM���xc��IP��@���Q^ur���� ol�3Ɵ���+�FF�/�$>aq�:���j�(a���[��Β+AWz���#�Sgk`J�;�e�ɬ��f�!��G���,~A�?�&v�c]J��p���	|�n��6h��bG+�ǰ<)���Z�C)���6L�<d�C����"�a�	`�����'yZ����]�g��Z�b2�7��A���Ǹ����G(�/�7�u�-�J��r��+�T���2Q/.��p���y��t~w�ʛl�N���D�P�7D'>�r?)F�O��c,�}V���-IԸ(q�X�#�b|`�+'����Z�ʍMN��Y<���S]��z��l�(����f�螢7A4���uH�^��;@w&�1#.�S����|%{�AEL�FC����R���R�~t���1ٶ3�qF��Kሔ����#�l�͏S���~B^u5�k
y5�[0�N��>�O�����RNd��提��R��c3}�bb��"��P�2�)
䨲ϼ�x{*�����m)�i���h���MX�����_�4)�;�=�܍⹫����"���Qn�@�Mԯp51t��JШ�-'�
�4+��`����к:��a�����ïLn�M!��sr�grF��v謀Ϯ�/�E_�$t:2g&x9A��"k�kЍF��G�3�VO�������w�Sn�&�U�U��-[��p�=�ƪ�k�k���,�wBd��5��ᦌ��
$ṗܑw�T�'Cf[J�㻉x2�%�w���C�tһVa�z҈��(^Z��clHPl³1?6и�]:�m�򮧮��6�X��( �w/�X_20}t�Ծ'�<$��,X�W�[8��t�8D��4��_E}j��g��sR�rh�� ����I.���@?�o�1�*�-u�U���0l2x�-�Q��4 tH�PXOHwj�J#܎^LϘ�;���z�U��A: ��(�<j����NB���>�jmT���}W�ô��LyPu�@dJ��c�h�3����t�e�*�R�!��H�Ѷ���~�l�k+@qK�SF�Y���������ǒɬ��}�|ᙱ,�G�P�ִ�;sN8�6�Й�l`�T��(�{ԐO����zj:���{�KZ��8�V4�i>1(gk��u�����M$N4٬����i��`�猅����)Q�:�'���ṇ��J�'S�,�� C�J'B��!�06b��/Ǝ��#�[5HQv��ڴ�O�*�o�� 0���'�n��3���Ѳ&�`�u��H=���#DGk�eX%�sʏ�v<bV�l���J�0�Ƚ�k��;m�NZ$*��Y� N�v�?��Ħf(2����W(��a��,BO���mdףo�(�ˬHE��d��H�"����FK�~����ZǼQ�i��,��HI�|���F�M_�!���~�>�J�
��ܔ܅��F���לE����4|��)�
�Y��b�o�w�����Cy�Ly����Ve]�G-��~:ɐ�}�6�����W׫�Þ�B��RҊ-\`�N|���vw
�*�8���J57:��ӷl����i��R%�0w\���Gա���p�d׈����*"]�$1x����1|m������=��[�<_���e�@���O\��m�Ϧ���������ս�`�ʲ������D�8yѺDS/׌vݲ���h���1��;�/5�{�2P�f�{�S�':t�Io'*#}�	�/����r1n]$>_ck�V�/K�B��lq��Ꮆ[����vP��d��R)�c�r��&����4�����!���5�jS���7k�u����#��ŷ(n!�[�3d�eCH�f��a>��g}dm���N�~J-����E��[|;�YqCѶ���)��X�W ����,���P@�.�D��p���\�K�6��.�>'������D�p��<���bׂC�$������h�0r~o ����ҙ�G8���(�	a$������3�UsM-^f���e���M?0�]�ɿз��T �jL��fL�{ʛ���=o��͖v��|�CpoŚ_e�[��������b襫!������:\�b�g6�4�5 �`�gԖ�x��Ų�"%9�?}���Q��T���dry����y!�X��	n��P�fA�(��0r�~7o����LKqP@�M�rI�����К[�H��M�g,+ �6C�/����'�Ǭќ�A��{�];+���:�mK�)đ��Z���a�N'4 V��L��OkH�7�<@�[#c�޽4�/	%�9M��*��m��X{�8���j���凌#�Y��Zr� ���ͽF8:h3{�M����%��Y�׶��c�8�茎�|@����
8X���S
�_r�rs��w��Jduٚ����nE���r��Р���s��f��Q�����9���]�g�\եVPU�5�u%�OFQ�*�L�1�d���ϗЮj�����WpJ���.���9���}���o�\(¶۵k�������f��n��#6�^N6>�3h4HP�9=���\3��z��&�0�x*}R*���Ƕ֮]m��C`��ACKtV_ɠc������t-������3�����z��$��q@!�C�*P�5A��I1��	g�B־l�j���.2)�Z���ewYX��oYkȍ��m�*_�l������9^�5Vq���f���h݅9k����TL9@��k�̿�cy�F�L���$�D`��DF/B��Ж�W���Ed��S:lR�ǐ%~~5X`��M[<?JؐE5D�� �0��W�X�>�)pU��YWV�-ָX���'F���M� �����pz�c"�pEr����g�o*�a�Tb���0�jM<*�����Ah��	����_�Pw&���kw��f��wk�`��߬�3�^�Y�� B�j�KTo�	˩Nf��UF!�r �Y�g���)W* �ډ����u�C�_5�;�ٗq�ٳe�r����a�G�~����`��1q	��k�~�f�@\妹�X�)�o��:r`d�5lTX�U�
�i�<=�����Gz�����k����	[��J@F��+��cȘ���?�ӭ������Y+�-��N,�Îq%��m-��G}��!6�?y�6�#
�i���x� ��s�=W�K���j-��&�0z�3.S��S��lSfh�4��t����ƚ���拉���&I?Åa{q�W򘁃�"����sX}��}h�U��E� ��WT~Z�����ɻ�&�u���\�-v��9#��Zm��ZU���#��W�J_�)�h$�g�C���F��L���`<b�A+O���j���9 �D)�Zp:���`��/�/��r�T��1�ǜu01R���]2}v*��<���;Wƭ�g�b�e�^LG�.X��THbK\N�1���������I�(9
��`�i��͗�ޠ_=�b���	��Cv����m;�MV	������'�/M�Y�f�� J��N��g봒/X��y�ܐ���QL���iѭ'(s�Fמ��'�52�Uf� ���H�����Z��.P
�Ms�#?�
Y����8��(@�<��]R�Ǒ�4N00_�$�ƛ{Iy�a?C���V.b�_��߉r��:�%�6ө�ۿ�^������ɰ-��8Ҕ�$[�?��#�/��<<����@�Q����#��<T.���p.Ư�!M�w�/��g_3{%�C�����F�Ģ���л:�9ޜIg��D�v���0���u��`s%��A��Qm%j���L�����ܞS`�c(Vg2@����_�&X/U;��=@Pd��;�{HJs������\m܏���O�u��(�/�'��	n�����L5r^>{-�����a���`2]��t�ՠ���yt�/����Q��
��!3�����w��-3���G�-��J�zT�
tG?�e֍�]�!��F+�
�=3���On�ץ�`��\����c]]Twy�'i$46�52�n��YE}(�@ȿy�f����k�~D#����i���x����96����̋&��Sx��%����e�:����a%���9�W(�˧���	cT��<���_��5��֍a���~P'j�,-��V���l�x �ǋ�cG�%���+!�DN�=����&��o��};�뼷��1�$�9�V�a�*mm�d;㯱 ��x��x�џ��;�kQ�z���"7[�����ϥ�p���Y�:����tę��e�O{�&|#����ו݅1�l䎬;�@��^�%����B#�K-1/�����:`����r=����0��ژ�x�ҳ�Oc�g�1��P/��z˩ij�ȹi�X�%�/g�F^�"k�� �X�a@��S�oz�i}�Ѽ|R�˔��	�J�s������ŁȤĘ Iu�ͩC�:���
��-�=K\����#�mJ�w�/�wD`5r�/ݳ�"T==~�ry���T>_��Bd��dT�@�۱�c~8K�4��@��~_5l�s�J=��1au>T�S�4��)�k�*T�E�����Jo0������Z�'�ۧSxu�����D�(�]��y偮/3�ǯ)w�.�BJ�0��<��C�Y�V��t�ܵ�s��W�H��.�pA���3,n�愠]V��M�P���� ��S�9�$�##�< ��f�8���\in�OW��a�ʳ�|vow��푒֚�&pq7e4�y����x��t��O�h�:�I�K��Ԍ&�z���sd�����aGs��	w��D�hk<tV�+�2�&p���U��Ά#��44M2<6�Tf*�Q�z���z�*כ����Z9�1�I��M�_I�{$��VK��t�G@��1��8��� M���^��I��
��f}
��_|u�<��jR����{2nK�ϩ~Iė�]}�	��v�ulq`��3��oҕ6�t�h�G�z�n͜�x��x�DL#����=L��ڧF�Ʋ/N��ā&ʺ�	�j�%/:���2A.K+~� ������)u3�B,2����t��cK�Op8��ZŶŴ�bb����,�hS��Ŀ�����z�2�"Vm�%�����%K[�!j_��nN��'�Q�N�������4��׬� S�����_8��\�"�f��V$�a�]Q�D�z�����R���<����:�ev;�ֵĎ�pS,i��C��;S�SپUVy��MN�2�D<�! ���sp���/;�0C H<��2�f�f��F�y��o�5j�<dE�"�/^�+W�y�x�y`}�f#��y���G� ΄�d�б�m�ʠU� ���mr�t5D,�*���u��Z��]*�^�J�,�~�@��0��_&���=�r��a����9}��̺��KRq�/FU�3��s������揇r,��a�j��N�=��WAM�ЁlYf���r�qJ��4Y��
U�2��T���$�l���yْu�XY������@��F�tN{��R��a9;FE.���*���i��)9���c����:I�H����i+n���yd��*N"G��/т/��H��Tx��1���@r+����.���"@��<hd�=Z��e�/�i�,� 8!Kj��E!� ���"�A1��?L��Uw"sVJE�tvO���{ʯ߱��a���p��wSP�L���r'a�n��2�`�|���txɍv_�V .i�n�n\zp%�7Q����!@`� ����=G0(FKs1?d���a�Gp<��-�ow��T-mO��Oa.WVQ��:ɍv��Q����m�L;���]y�,I�Ǻ(��h[��0j��C��y.��(����f�x��\���Vn7汢����fF8`i����t;i��}(2~��ޭF{���	<*n��'�n�ؚS�!ٍBQaބ�Psjy@߿:�`^�8M!���\��)V�Q��!���/�@�h�݁�|�I��vd�� ��]���LJ2L�馾��+�'�w�@�v�Y���N�VٺN�8_�����uՏI_�iPZ�_��B�}�g��2�S](\FxC@`�	�a&�޽V����}���7��Y�S��>��̿	��gZnV�C����c����B�@���cH�_t�c��QO�[|]<;H���A�'��2�\�PU�9���[S�$��c�T	��K��&'Q�D���c���36 ���Q�n�5����^z�>]�C��BC�l����;{�@2J*j%3�_�N܋$-�!q�	��cIN ;�r����	�E�_ڵ�j����åE0����0k*����c�䏑'�؋�f`HӷcL4���M��oW��$���w��8�6���SfXC�$��ݓ�E�^��Z�s$�Զ�:��0S ��[�{�%jGt�Z���I'��]b��9�R�d��È�kr�|���h�7� ��H��8z�����->��-�Z�|���̓��4CFdǾހ��C��l��ڢD��ϮMi�|Ǿ�>X�a�%���/lߋ~��x���=>� �z(�.c����?4��t�Řa�I:t|
�H���^�]V.��# 戮�.���q��M�
���{�s���1�`��oې��� rݰ�_�Sum�D�ұݎ�m��,�m*Z�����'�L����	Vs�ɂ9��Mw�����<���2Fi���^	����Ca}X@�q
iǒK�<�~t�����A<�9V�^3�]P{)ٻ��=�\Qa+����4Cյ��/���$g�{:�b15� �mQL&�Pg+6�'q�0L��VB�s���w?Ӻ�
9r�ţ�#j �0�$=z
g�xr���|#�p}S�/*��/��5�w�YL�9Z��	L���̮A�>E��F�bAk|Sb��4 ��l;�Ph�j*�u���K�!���I/�$a3�\L��1�H�eL��Jv4@�ͳ�;G	�Uծ�(�6�M��8��?��h�n����[�H�@R��Hi��kp��>����2xB�t���
ör��D��nL9�G5������zì5�o�v���L���B�:꙳�P�ɮVN��E��F|9�9��oq��ԧVI�o�=d�
�ߔ��~�1�4<L)K�Q�P$��Z�ڦ��eA��>,2��Z1ݭٜ;csK)�+ߗPwF-�)L�q	�/K��5����FQL_�5D `���Cl+�`��c}�ݢ����N鏷Oqh��9��P���KC22�U������1���J�D�tѦ�+M�QL�����%����� �}�g,?�����65f��U2wf�Ż�3���]㰿c�5��nI��Ca��D)�4@Ύ�t���W:gS�Q|������wkx1�W>�kR�b\Fd��!��7�Ss�{�p&kk�{�p����Q�S�ʗrv��� #���K�y��[�K��7]���y�0�����%Bqq!t�ު���!�< dh���9��LTh���$�E��Ĝ���e��4;����um9��Br���A���;�w��K� G�Ed�6�,�'m%BҶ��S?����Z|����p���T�� ��U�d4�5U��%~6ff����\���4��s�{}	_>^�,-Ɗ��z(j��Pp�v��|���g�L�dm�6TX�qW�������Ags	V���D�'�Fm��|��}y��� `�j��D(J�/�h|�b�M&*2r�ҹ?5!���g��]���{3c��ק_��^ѽ�Fq�Ssa��Js��
(ua:¾���cbg1�CDP��ٔ�}l
?��y�]��(��O���i��)�?7��&����WL��iL��t�y�%��y��F��hg:���?�0V{��id��]:_V/�>��rݸ"4.�~�����ֵ�{��-��	)Z�&�z�Y���>��{�<~@��g�k���Fk�eH莌�i���,\ѩ�V߉L�D���3L�0��H�~ښ����k�X�hX \$��^���BX��N즢�P`�"�����"�ԟ��L�]���N(�p�Pa�Iɩxȟ�r}�b�uخ���l��VP��u�Ԗ{�"��.TC&*�8��<�C�	�M��xk8i�$�Ćr2C�=�A?�H������Q����H۹��g������l�sᱍ�.�n�6��?��ys���\�N)m�nPs���U@�[jF�x���Y�ۏ��:N̠�_I�� ^���l�Dp�p쁑+�������jF�)�<��)M�oR�D�ÿ�n�!����t���99����7��~F�/��X�Vf�غ��B^�ڈ�h~����}Z��
���7���C�RNoaSh�D�Z=�a�^����Hs+|�wǬ��ۧd�9>|�q�o�C����L��wư^�}v�g����ߢV
�
�[�DӰ��^/ҟ4,P���=�_�3b_'9��-�a���[���Yp8Meu*��f������:�pfA�ʝ�J�f��>ڂu���ŵ�����(�Ft�H�P�,�飽��_|=g�G*t����ԅ�yG��j� !���P}?����A�DL�1W��=�� ��"w����m����m�	����C�E��n�,�������Ce�����Mf� �;���WJ��A��7[��"�b��K�p�M� &w��ik޾īv�E��7Z!��ږ@Eˍ�:�	����v�)V�LHfȆrp0�a��s"77C�qZ#�o��Ҏ���ς���.r�����$�5�:�ŀx��Di���I���i����
��6`!ȟ�*sٻ�x��;N�R%LyN���Jv�0'�Ѵ����ZY��f-!�T�8��Ȃ�G_H�5�q�A��}�k�v�NZ�\=8���]۱������K�:�Һ^M(��@.b�\��M��Y�WPp��)d�|�G�"�7�0���9v{`'I����j��|%��L%/w{(�`%���������0�;��pϔ�a&�T�)�`P^{�<������P��6#*9�YR��(\��JJL��9��'x�sϽ��'g	*�ʍN$��c��*g����Y 2P���bB�1�D����DY��IR+X��#�;l|����ε�ue����~�š���p�b��WC���6�Ÿ�φǤ������Z�Ż{C�Ɇ��Дx��Iq�����dW���}�;`t+��[�ܦ������F�$A���"v�5�5"�
��xI�����Ǯ.���G�R�%�|��h���iQ꘰&�g�?����X+5~���tV���e��X*h�Q&�߸�vC�x@��4�E/�ڐ^���[q���?�1�B�&�����밞$f7��ZĘ7�Y���}�:���֟��ӝ�I��s5ɿ�:o��0�Ǒ��#w�_�?��W�o��$r�<�67����P��	?�u�L#��~U{�F��jx�WB:���/Q�a�#��/���5z7���\��ڽ
�c�|���������������4
�i�q�T3�6
�\�I�:0��"$�(�=�n�jI6h�'��� ��>H�����1��8U���,̧�I�-�Ft��~��T��p#�3�=��P#�|�=H��3������^d?*�ȶ�/!����`�h��EB4��;�>��L�{c�{wu}�-6��'�7�p	�Q�R�R�rH��,�F�Nn<�t�5{���dR������'�k�T"ѱw��4��Ii2C�[��ޅ��B���M�|D`�V�6^,Z���G���\9�k�k>f`?L�y�c��hI��^F�R��cJ]�+ٷM��W 4��u�4p��|��{��p8�*+i�{j���+�-w׌1��5����In|��9kGQ��c5
���,�]�nC��W�|�_)��BU^�:n3I(.��*�g�0̆�=�{���$����p��zs�o������x���2�2�r\g@i��f2N�zPWP� h+٘��sWӉ*�!�tbw���G�n	WϿ�R�����g��:�.m��/	Ũ��(�a&�[ r�CT'��e��A�8�����4�����|/�>�i���c�N:6�Ir�Ư��D����B� ��ѧ�׮�R�hW��꼶���/UMvo��,i��y��@�@4�ɴ�nN{�)��J���/�<�:*��	�!� (�ٗ6��0
*|Ֆ��7��R)�	N�/N��$�q���'1�;�[��=g��i�Ų��Ýo�5-<x�����d!&�A������������޳c�.u%#M	ӰHM��z	�|)�_C�ua�m�f��qC]D�:h����8�.	���lt���٠��oh��7c�Y;�^\���[��-��6YPX�6����Q�����Nwa��f�����q�b��q3�`+q̺|��yHl(��[
B�����E}W��e�gúJ�:�_��co�b�u�;Тoݿ�r)����Cu��;=����o��7��;*΀�Rc�&G����y7<��u;x�i�4��c-V��-U��
�;(BF�w�IR#t%����
7���F�E�B�8�ÆN_�s�ɶ�a���#m<��Ⱥ��/�1�ҲI�=O�x�}G��
�-`SPV�aEU���lo���+P�`q����
D�ƭ�͢�M�GmJ��i�j�:m�ʶB�6�pA��O3��
A�U��^V���C�p�:7ĺ�=V�:�V�RV)�Z���K��@��^ڽV��]]"k�S��O>�V�0��6|�Rg;�EEpf����K��ZVXJ��lB���6��R�2ǒӾ{���	��N%C�SwcI�Z�A�~zW a�z��@���_�Oqij=TY��.�Z��#=q� 	�e�����Ѩ�a�LW�?�u�r�׺�8q&�p� &�Dt�9�j�1�{?1,�Nr�K:�6�_g!4��1�Y��-p��7�`���^Z�Q�ݪ�z� ����UǑ�����qlZ�A����C0,�����N̰&����P���9a��iRV�N��8��d�Z`�ʪ	^*�a�w��菎t�R'��	�ɫXg�wu9=�,�%��[p³������͐ÿɗ�@�OjY�z��
#y�s����TvV򏚕�
Ҷ�����e=QXZ�����C�؀��	�_�YlT�G�_��˩`��e�� �㩚q�UW#��*o���JI�n�qd��"�S�3�F~����tuB�G���G>���s��$�q��{\�s��� ¨԰�ű��`-a_{�&1�f:�W.���H=�r���)��u�u�ۓ��|u��q���(6joW��a���E]l�Gq#��X�>c�n?��-�\���S�;�d�{?yc�b�~x�(�	�j�&S�h̹� ߴ�u�x���/�O��z9A��kXZ$���O:IȞ���R�E�f�4�^���]��,����r�$��~�=�h^m��B»ooɏm������*������o�+ F�N���6K�& 6���������1X���K�$���,�<$�d��Fd���`��W$�{��ϏmTA����a�L�@��=��R��E9@�,��܄_c�
:]��p�)�?ȷ	��"���'Sx����9�)k�O�<���8�睈DX{�V����}�`�P,��i᫫x�5^�u���f���~W 6�Y�e�>�Q��I���'��y�iĺ�u3Pa)���Y1�qc�&ҩ�H��PdZ&c���\���JL��!6���>k��e����V�I�w��(D�|1�JZXb����Ʒ� ���X<l�����^P�n(N�g��cǲ�()*p�>���ȩF�����9��U��������4�K��Gi5�(��6ֳ��7}:4����w���V~�=�m��由�#5VN CRpt���H_@4s�s;dI4�u�y\�+h��?��c�����lR��J����&V�EI��J2tU����d��V�5�9(f�IĴ��vJā�OU:�����ђ|DA&�]m:���@:��o�t>�5���*t�tj��(z@�q�pi�W�Ud�A1���Ff�ڄ�����yCc%�)�Dh�OC:|���;��Y�.�D��U����s�^{���AIS�5��r�{�����TX�u�c�K�n�"wI	b��%%tmsaW{@H�Hˉ�-�R����lR��JL8 �F4Y��m�:����s�f�YB�����x����|��9��%q84fp�2�!��\���1 �`S~l#B�z�79q4r�%�/������E/������v��,�{���=,arK8_�������9��]�E6M��#�M�p��p�^� ��J&�ri��YiW��L��d��=r��3�+0N�)ƴ��F�>:^�i�I�,������j3AO��]x y��j+RH�b���jKA�q�P��c�.3�d�#;��B�_���>n{�-���R�JD��i�6.�IS�c��
�=�;��D�[zC���U���*nC�ذ�8UW�/H��Ǚ�%����m,�#�A|<L�]<���%��JXSd��*�q?�K���8�z�)V�bmQ�����0#�f�c#D��tdf�����0>&��Bw�uM��}z���lT�%��J!���j��zZ��p�&�?44�6�Z"���}g�aV�����f_��_��E���1��B\t��4�gV�Y#]�1^�7��),o�\uC���1�X�C���x'�'��$��I�莸����@�:Ay��Ǎ	�(��rv����O���ժ�L�K�B�#;7VYw~�[���-\��lc���?\�N�2�<UJ��W���J�^ki��gc�W!��1�$zC����of9����������r�8)��zW�s�K��;���uJ�-�ʧzN����>��b-�Z����h��T襱�v�	1�*o�:߻dz?��k�-1?�{��~1�{<��^�������o�}dBC�l� ~G�AE$��&��|{��</X�)��T-�y�-i�)U���!������=$m-�hm�~
ދ@�/�`	�o�4�����N��(��S�a B��rD���}��n{�A8�*�&��!%��qiڰr_sN�,��Ԃ������22YR��(�Ѕuգ�U��{�r�u�:8s¢����zyz�Y7D�ڇ��پ�3ȑ���P���G����$�B�gP�S�aⷲ������f�߆jx���N�I�w�Ặ�RDԜ*ȳ_�rHo���b�s�{�:O��ԣ�O�/ޙ�*)�k��D�#��M��`��j�M�@��ǜ¯��R;b/���2�7j������"h��dDE\n�ChY+.:�'#�	$T��<�T������Q���{��;?���f�/y�����U�G<�rP7Oͯ���ǜ�Ow��ƚ�����ĭ@���]B�iIwΩ=��l����&�5�1h�g-g^�J��v��l�^'�!J��p�����N��/��c���L��q[�_�`�@�0���'��A�+�'!�E�f���޶��Zqy��
����,�F"���3���]Ή?9����M-2A5�ER���S�2g	OG`BSM��� ����+��79��3�S`(N�ӭ�8�&gv������
y@9q�r(�&־/�������[=�&�m�ڤ<���Ռµ������k�>Cg����$T����ެ�D<��!:�)M�$��:�3�1�j���(�WhB��}�[��U��R�x!����I7 ���0�@��4次oWЌ��~��6�G��c�f�G���硈$d��u��r��}]Rq���ĔW[���$������{�\(�S��T���6  ��d^,w.�H�h
ƀC蛯�J���ZҺ�
x�L:���1�. J��$��է�#�ؒ�J6֪����a.	��Qba�s5���vY���Ćc� xx��0�߈.��ap��4G��p�%���d@�_�1�����F�?�*��Ԍ�V���'�Y�h�p�y�?��g!�?Wh�\΢��T'���`�Q\�!��ϟ�3�>�p��V9����Ux�_�G�&�+�D4S�0�婚��x�#$�f|�k)s#EPD#�$Aa閪aI�Y%TÆ�{�")"Y��x*�L�ӿG�TMB ���VyIE�5���>�M;<��|�RQ�.	iu1�@��̢=�Gm�.��������("� *����jO�Pδ���|��6�����ҋ���8μ�5�#!!@Z���r������E?�}ej��r�@�dA�!���0�xG��yȼ�7�;Q�b4���1^���k���$sE|��T�r+�l)���r>���3���� �>D�v��ɔ9�`1+9�-��?|p������o�k0f�@�.�"�_2���bQ,|]�S�������
|JT�^����o���-w��֪	�)ڦ�.�ka�JO�mG�zӝL��d�|Jю'F
9�#���Z�� �
��fU�}s�n�30�V�����m2�7��X�+7��o�V.*�
�ڳ��{f�f��������ڴ�>�Ƌ�J?�Mz�Y�z���':���(A���� ���p����x����3<8[#H� ���#֚��y�L�b:��z�b��D/�9�yg�)�� ���i!m�5�e�0��T�E��߃��>%?�;�]3h63�`��q�`��X�A!����1�XH^T�1��`����^����i��nR���!�e�1S�]�"�!Yk������SA��w��Ȣ�ѵ�}�z��J��,��?�R|��U%`O{�_x��<!3A�n�:��?�jw���'�kJU�A����s���s�6�z1�B�<��7c+U0�=��
h�xc͟Rl���o�}�d-XYd���B�q�H�c��UM�)��؎�
�_@�D�pUx�U#q*Du+MA��.�G�Ε����(����`s )T}��F��t�c)��%���T7�
{?�d�c���H�t$Y��Įa��23��Ν^3r'�%�+A��ӗL�*p<�����I �>���?�Ĉ&JH�+�fI��4k����0Q-���P�����|�B�
KV@�|A�5�xA!���1���MS]�xU��6#O��g�EDN�JNx���Q~��;��9#��͏{��c��P���j8q_z�B����.墮��3<ʔ�ipY$�,���>�m�u8dG�Gio�V����� ��Ő��_����q�L�)�RyGQJ� ~MA�l�|�?�~Lˮz��>���Q��2E�X���b���7 �:�&W49�@t�������,�F�p���	v �;�������R�5���1�y���>?<���p��jia�BC6���U��Xw���lt�x�����s�Y�a�C�K�[-B��,h�"��?	�ev�F��z8�:h.:!�� �v�����g�Ρ򑃔���Z��bq�vγ�6a��jl
�R�1G�w�4],�{ښfm��6���%�nG��UcZ+���r.���Ў�,�5��a��Р��T1�x��Ą��������X���fOVӹ<e���f�P���'�[ꇵ�IY=���9���ʣ?���"c���QZ*[VƗ]ɗx�`e�L؟&V}ʫL��5��vm�.]y��1�yq�+� ]�&*��c������y��v 
9�_!g�~l��"�A#��Z����3�����0���ٱ��z\�BD	�lY:M�f2G�Rh��a$~_
H�a�I�s^:M�(<ڣ����mj'2�����
���!O�afN�M�i�N]ňʀ��a��O\��m�z�F
��n�g>D�h�Sp[�y��n�����-�@����dnΕ�,��������
͞���v�oO���w�0@��5�V���ߨj�`N��u����X��h���'������\� �zWcp�K7��fV����}Z�C]Q� /�kӗ-Z��"����/�h�9�<�T�{�wB���
��l���b��ߡ���jK����ۊ��"Ս(����GZ�ҙ\��^��d�K9TNٷ.>x���_*�k�t������/�z�T��p�
�����a*�}��(>D��;j����^o��&@D{
B�쁯Lw���zTj@)*`����	hϲ�ك�D�Ey�ڕP���^CJ�7�M�|J�UtWR�������u�?����V^1�Duͺw�8H�0
�u��Wyȫܴ2~p����HX�����v�¤������}V�g��%��������%���L%���7��d��������%Ve�{� ��;~�]�`��Y�:���2��U��I�<����X�_������3.��]�}u,�|��j�b�21�K�b�<�r��<g�6Sz�����G�±�:U�`��#�|ŚA%Q��^˜�-�C߈$�\&�ƣ�
Z�}��g�b�>��`�s9��(%�c�����V���Jѻ3_�}��1��<`~�N{���BǾ0ƾ�s-R�p�@rx��22���+J��c�|e@��-��*����4Ѳ�y���F;t���`>7�[^�|�'���!j�$t�+��\��ZPӪ�"9�RΣl��#�&}Ԕ��tsr���W	���j[�"uZ�j�}�w��IY<��-�t�li��9V�)��n��_��`�n�3&��>����|�Y�*`�z`�zZ��8�؟	���I���h��ԣ�[1Ѫ��[+׼���A��p"]�f��Q�SƘ�AK��ά�4�0=-�k����Z�(�sX�����mK�bX�l��rq��br��L�#r#��U~���[��fi0�1�o+i��G|DL�a��;���'��n$���}V�b=�0]4<Ѿ���WA/<#�P!��>l�O.%�Uj��:z�Ǹ~�P�3/�l���O�8M�[\��X΅��N,oz#v�4��C���Ŵ��[�v�]�oV�>�̍K{��&�]����Q�c�B�|ƫ�p�{��r ����E�<[�{���}ڰ�(���g��e�߮Orȡ1�>�;: �<K��^�Ay���dd&��%>.���|��{
rGP�N��7A�� �8iޕ��B��d���2�f��ְ��w�ӕX!4�#��e�a[�����b�>���=��6�	4JK����af�Ӑ��T�$�(��K���+���F����G���iT��%��q�f�×{<��k��gx+㈼�\a|\���x�i&�������5���;��6:>u;gU�N��Y�A+#�Τ�kVnÀ*�����) ��,�<�)�8e4�^|q�>}���{R��^.)C��ׂ��6�Q(]�Jľ��8Od�_?�D\.�Z�;G�V(ޱ`i<v�4S��B�҃f���$Dj��d����6G%��&��+�H����}FwFh�ot�g��Ru�Ƨ��u����*~�l�JR���aJ�ϛF�9N�y��p�NG6�-�?&��=-E�
�R_�%�?����}��9�Y'0f�-�l>|'A����.1ث�:O���5�t�Z[S�yA$��2]�1:К�X��ϋq'.�x�P"ep�~���qn!i�u��Đ2p���` f��f�������,-�-a�h������v�@mq�_���O��QdQ�}�飳�K�]l�q�>���B\^�DfN�����§xƪ�*��$�Tê�4�@��Fz넣{/7|m6
5)�&�� �؁P�w�����M��q�M�j��Dw������)�Rb���=��-�R�R%�
9{\vG�H��%���`^�[\]R,�Z���(����QC�r;qM}.����R��j�J!4�J1f} �91v.j�f�Ё����MM>J�pƹ�s��~�\I��x4B=6���Z���08sejfYTQ�ƕT�w��̬��_���w���-=i�H��<�s�=�g���v�3��o
9�l$"��w��DXf]��S��
ȯ�jX��Kz������I��� n�r�,���fځ/E>�݁h��ƀ�|z`^��ѲjB׀��rts�]�G�B��4&�!&2�4����� ���32�s*��pFX��(�itR�E�\��@�6k����S�O�d.h�vx�>_ϋG�[���`#B���Ie*������`o��c¢jho�m�{��ֈ���S�⛦�k�T⋲�c��&BϽ�q��{��Bx�=ΟF�o�7�q|�Ojv�������� ��t��28��2X�ȧ�_�y��8A$ĸp7�����_l� A��"\{y b[�27<�	�l젾�Ĥ�lT�d��uc��ł_A�X�c�(vG�"�o�f�b{w2��d�a���W�$pIvb���t�9�
<��=��MC~\�f�c%�Ȣ�r�c� |��Pͯ��"Hp�|�������g�=�6�s��f��6I��ڄ^�����-���T�|��1���<~�.67{Wi��uY}��	SldŒ�< Z��5�Rk�x}�<��w�����N����dK���89e������I�����N7�UVg��x'�=�S��.L)f��Ø�[�2���q�Ÿ$�SYL٫�˶���	���>ě8F �4�ź��U��d��u[l	0���}�s�\��<r���ҳ/t�֝�u�YZ���A8,?�T�j���k����=ʁ{<�$�P` 8W|�C�f6�̴�r˄|3$��o��f�p>�Rx��7qQ �=T#�Q���sv�x5"9E������p��b>7^}���B���[H_Ǯ�3���]��ׯkb�T
x�8ITem�Ĕ�&�]^&e�X6��B�Fuq��GΤǎη�
79�Hfy&!�j3�P�!
�N2�����2�����ow�ߗ�쁻��eL3b�!�1h�����)_��D^/���q��9\����)���:��,j��b�L~#�1.���ϊғ*��[���خ�l�����>i3��p���n'�O��q ㋁�?@ݮRչ�/ݙ�`(���l �<^�K�}WGħ�NJ�h�A���˷|�۝M�Dܢ�"��iB�����$#)H���	�4tͰ��d����%*une3[]�ь��h&��cY��z��pS`��l}BYC6����g�����g;���@�ӗ�5~+?�` ��e;&�T���q�^4q�V7�
C� �(!�`��¼P&�_q����~o���'�ʻ�X�wu$ei��A'�;��=tq}�1���Gg�HVqr(��<�+�e��mg��r�)\�}¸���$���]QZc�ۻ������+�KݎT�5��2��M�L1�rv� MҔD�l�q�8�:2NZ�x�*���e�:0Ǿ.AUQp~�r>c�xZ>2�0�Ϋ~��r������#�/� V�>(�\!��]n�s��^@L��ZHZ���M����Rep��2	c	=�o}�����8��*�\ٜ���n��@�|t�-�'�s҈�
o��@��	$����1�"���5���a
�!78V��ʫQD�%��R���v�4ם.:R 4�!���ŕv>�{�{U��R��f`J�C���fqt��N�4<嫭�9��]$h������@:s7��VD\"E�i�n�E��,�s@4�̚�d�7[mo��u�����J������qNio���޳���?�m+N��j i�^����2���I�7���\�V�d^����n��J=?��T1 ��Хa�J����׷��䁗��NԐ���9z�wd���Zd�£dG��I)��Vfy����Xz��-j呔6�,p���&`EZ�h��H%j��c�"�m{��s�33���o����T���D�uކ��^��Gi���T�����>�ws��<�Vmn�[N�A$�HE6/~�D�`��l�@%e���jH%=�*���4E.�L�hB�򦬦�hl>$�]8�p��6��4������>�@��QZ�@��ذq�&J["W7)��;4jcƈ�O1熑�D �<�������ɏ�����J�����.�8tҤ���J$TH
79�v2nTJ�0-^=<��`v?"{e<ƝC�ͭ
y0�I ڄ��5�1�G	����*�*�=�2���7fW��w��k"���Q��PЁY�ypMbi�A��mnl�͔ �T\#O�Z���ɯٴ�����k(��0mp?�p>&�]�t��f��T����!S�)���;�;-�*^����?DB�;�TؖV��`�?Ge��4��狽m�.[9a�Y6H(�(��*� �ʁ&�[����n٪p���oG^�$���Z{�u7I����7�0��}(�O����T��}�l�?�n��O���������
��'��x$}j.z ����P5)t�+�{���;�q�h�QH���Ö�VJ��W�]D�w���v�E�s�D���m��ZK%2Biφ�ӈQ�&���Y��I��C��d���@���Q�uc���Y�)�6>�"-���WOl��2����?�����fJ�1|��r-�w�dC�'܁Uj;���R��#12ҿ�=2m�t[4�e���������	U*����A��e�İ'\F�m>x��F>�b*7 j�}���F-�rP2���-Hb'�*'��q�p{@ٯx�~]���t���	:a����Z�������3�*q��_��`'�Z�:�0[��#e�:K�S8Vm�J|�HE ���S>$[�0F��v(�׷����O���U0��>��C���; k+k�>ǟL�)����K��ýt X@�l���k�x�M
���a��)W�k�����i�On^�^	�ع*�񷲑[�yɸ��Ԉ'1�m�Ք�#e�Ϗ����kA�r�b���ڻ�$��)�GY�N�6c%�¢Z�ZA@�S�qR���U2���H�lwANB��Fd3O �w槞�M����Y��!ǣ�N�ҳ[7B�m�LVE�K��o�T ��w2N7M)�PLM#�!�C�E�k�<
y��#��VRL�y�3��q��|�4?2�X��7���$��5W1�E�즰5��$<	w朇e��n��B7�s��9��j�Kv7H$̊���&yb�dv��NE�����ۦ��������UjA�	�.�U,�"���ǜ�)ܷ�^�N�7��e�(��8�9X�f�L~X%�%�3��6�==��)1��(�X�f�����V��4��c�E	�����.7�z�֝g4��v����۹$�I7_œQ`	�HGZE����)
o�p�,�/�g~�����FET���C��;5W�&�Ld7)��S��b��lF*t:�����gmػ����I"�-�o��򾩫�^ YI�2`
Ǆ��-6(��dOߞ�'��΄IK�6�P�e�]IF� o�������eZ͏���nn�+�n;���b���l�ۇ�+�G qB�@LdJ�wx�U�����?4R����0mO����L� 4 EA{����IѶ�sgFhT���B���,�]�Y���|�fh���D�"wZn<;U[���rK�����B�ԮW�O��_Y���4�����$V�B�@�����Vu�{�׭\��m��Z?�9���a�]k��'#��|4ɋV��χ���xV��8�]v��lÇ֜'�u]P1E�:�1A��Mu�e�q��&��[=lw]ͺW���^��CA5�q/��n���R���:
��^�`�c�7��E�sP,�a	�AG���X�
ƑVg�� -)�۲�����'�;]�n�_k���Z'@��) ϐ/�=[R�N�FxŨ�>r<�Cb�,ZVŨX�Q�g�a�>�5�4鹤���r!኱�D}I �M���;A3��=*�d�J:�	�Y�N�'i�8��ҽ�p݂�hC��� ���Xo��Xf��2GN��n���!줂����C]�����>��?9�Ї�ý��ծG2Kx��m- *�wO�$����%�������k��!����x�����0)*��*h)�c�^����D{�w~���o��ؐptv��ZuxG ���$�n�!�Қl�w��	��h�]�l�c�	XI���;S���d���+K�����_?maQ�c��l�Ҁ�$*����U�+����U�p����1<�i�<o����3������A�ڽԉ?�=�Q�=�8������(��v���~oN�w�_�z�����B�����Pj,��y
��] �)�݉�hK<M�z3C7+yA��5`�q�[�Ǹ_ǵ*0��뾐�%l��o��I���"�HNG�6�}���x�j~4$�%�F�?��-8��	���N3��e� �$�3�'ΛR\��,��l�	T ��}��㩉~�@Ĝ~�Z�DecW�ğT�)���M�k�M!BM,�"�s�l���F̖k��W7D睍�Qj����T����?��7���>�ڙ�ŢdH&i/����0VU�zV.U�MJ���Y���Q>h�bg;�#[i�7p/�A��@}.}�
�\o�^�%WR�@:�Q��}�����Üc���an�T�����7[����ބ������A;$�ʍ��q��l����M�P��U��D�9C�a�7�y��@b�-`�&���Eܼs�J�����m�� )=�G��?�{̊�v�-%p�Uɉ����-iW�T�`Lf+��)b�"����[�Ļ+��.J�'�bH������uߐD��������d ĵC(g�LYp���﵅>��l|��-��^�J7�}��P�u�)�K !SxSQ����J^�w��%-��VY��%�d��x!���+bH0+hX� ���Q�,��r�ڭ�����mr��<iM8̭IEq�$�N�T� :�#	z��5?*Oi t�<�D��K�z_�xg,��uKXܘ̻���tГك�R������6�F����S���(A6��;��R��ے��,��b/��	�<��L���j߻�Fk��"�ɍ��t��|%�#mI��|o��SJ������u��"����%@������6�@9�y���M�9�d��Z�ۑ��E�9�<�2���&\,v�ˋ+YV�����tZ����2��o��Y!�%	*��G���!��~�ā����b��D�9���܆V!��z�{�D����Gt����#-}�2�Z��Uĉ|�98�ZVν@T�������E��WK�v��V��!����~��e����CY��F/��_/瘕Y�d3��WC���21+l�~J�	������z6K�xq[�����$Wu� yd�@Q��E��9s�|5�3Ќ��X*�_S.��5E�0��Ձ�e��ꩭ��a#�ھ�@��]n1A��\�l����p�o�
�_3����4�����?����'�:��.��ޑ�H����:�����R���X���݁�� �sI�����s8zB�}�vā��:صΒΔ�e��r�"�ë�etC�5�7���2�`��P�+ܿ3�ņ�㑍­P��ڦ��_�[۔o���ª���Z.P�� ��-LG��q�A� ��V��l����#�7<�{U8��9bh5n��|J������BzPW]N=��o��Xys@v�؉�[��{>�Aa>!�~���ZBC�K[?Z��[�����e�z��ej�������p���%ŏ��G��sH��^�"�9-��H�(-EY�Tω�/6C6G��U��n�"}�4��@q��'}X�<xF��Q��~��پ��حbf�U���k��R����u��{ �g@%�"ZM��7W�o�i��.��k���>�P��!�������R��?2��9��l���l)F��A��z%*��<�0��S������r&X�&P@O?�u�f0��?'uVQ�"�GRu�
"�Ǒ�${߽U��V�2��=��%tÅ��ƨd���)�!�f���T{zR��R:�N�R�'���7U�ɋ��f0-���o�ܤ�����n�s�I�7���d>t�� �����$�!tI�i���I��SlW�D��
 r�g7�wruULv���g���rLD�6��U�}���㡒�K{:S��xJ��2�o��z�+W���b"(&�I������"�O�St�I�M����u��5��l���&~�eOF$��[��ƚ��;��8�ըK���R�w|%���$^ �Rq6��A��Ad���2�BRЅ�z`�.NDs�8 �Hû�j�M��F�xs`J�{I�����mpҹ ���� ��܆�g�V�,�K&L�j9�ȶ��}��������I۬�������*�CE��k�[�P��`��GQ�>a=�fn0I��_+mBk�O/�%z�'I�܀.�'�elY e.��-W�>cS��E1��"P���y�����.\N��*��WsU�~t���F�w|�`�,񃕺f�j1�u��4M���+�̟7��H��a� <���
�Q�`J��E�mc���`�K�*�Z�V�p��_�G����m�H�p�������0�ϣ��2
��bW}R��Z&�]�;9Q�EG���\���*��{vf� �C$�<T�y�z��:r�չ�嶐�!}��U֜�@+u�3"�S3��Л�@Zl�Qnѩ��E�H��n(�.F�)}���>�����ob�w�1��Bê�H
tx����y��}�.�+�DA�G/&�1�r\E���NƗvة(!�P�c�y=���gS+����N	^`�(q�U����ݪF�y�]�kFy���ñ$�َdEHqā�B>��u�\� ��Y+I��"r0��)��.jꣳ7P�ކ�����V���'�f9[^%�����4Bsg���^��.�P'����]�Q��x�![���.L���E�%փ��a�|9.?�k�̼C�c��0�=��n��]c��J W��Vzį���ʘ����kH7��jQ��a����U�z�p�����ps�c�RSP�s�|��O?��F��ka]T�Ә/��zg��[˛���*���q)�W�/ixMn�Eo��ݎ�P<IwW�x�-����Ǘ�F��~�.b����e�g�e�+�s�\զ��ǮI�±��EE�yړp'�gu�7�Bz�ȝ�O�q����� �(+��r!*i>�קW�Мa�޴�c�d��D��7�7��B}^[���7�=������+x��
��ڳ�g�����ꔛ??Z�E��g��Em�i�������� ����'�l�DczX>X�~�	"�]TkU�/�ik�x�FBh��Co�j�4�+���ML��Ϻ���T��/{^:��}`w��*Z��w�p����+n�TE"Lp���}�D�$�vk����3QgJ~μ��hm'��J_TNy��j=��{D�<M?�Ybǒ7�X�dN~B��+tq��U>bl��8��	&[&@Um}�� ���9b�H���f�o�w/Y�7��J���K�+��8�Mt�ZM������Pm�䝥Ct�ڲ�vNi"��q�1"`f�ϭ/ŀ,}�_ou�(��H����?�>�?��Ip%ؼ�0��9}��;���@�^�|@�70�L|�e�s�Z���Ў@s]�����H{����>߮��$�[᭬�h�"O,�����0G����A�.�"8Y������⌈��)a���vx��-�1�^?�ٲ�|�k|�aă���[��@���#�-&L���y��?�}�=�1�g��'�˧}��:mT4�]�G��F�mŪ~�@�ş!��D�ׯ�pC\�Eo�O5������c���hQ�9��3d�<:ؕ��#��f����*�Ȁyפqu��CYp���$�0;�v;���܅�)-D�z���	�SLN����)���a:��~%6S�2{W^�s�F��\Cj:m���eč��g��I�x��Tl��T��;䔼n���>�q��,A2��vb�3y��{�#��O�+�C������d���Ň�ł�����,#F�E�����Cd}Z�FH��kDzx�tvU\'�M��p����W��t�P-�v-��:DDM/��3�<��'Rs��3a>��/:S��/�T�K�6�g�=XF{X˷
;���#������T'Z)-ِ���>����gg-�l�4���Ÿ�����x�q�hhú� j��� {=��٪a58���FB�ww�>AMV��`ݥ�,��p8,��F)(r���=�U_k�.�S=(�����Jo?ɱ��hP���b �EYÃ���ʘQ�*�f
��e׿>R��x?.<�>2l٩� �X�H�� �̦p^W�ቺG)�T�D�v��B���l�0�m� C�Flk��ɴ���W��5����x��B%uiȥ�C*A�?�,��B�q��Q B�������dE�j�6�G��_�15HXٙ�Fu=��i8�;�u;��N�h�h���z���E_
�H"d��x��5f����j�u�q� ��oC����[*��&��R遟���[�u�^@L����mf����,N�i�C̤oE��O�[`"\(�t�Jp�xM��b�ws.�|d���{P{��|NY7IĚ�^K2�T��}�x�0H�q&�+,�F��U�K/3F��N�)m���kK�s��.{O� L��n�;ۋ���aFy�!M��4C���⌭ �Cni�R�7�M����^f�� ���`��� ��b�%�a�� Ms�
A�i���>݄+8R4�*
#ǒ��T_�&�R-�-)���_��[��L����t׿h�}�w<�2�v��zt��x��%�	��^����Ë����M�>.39���	:~��>������f%��dHfKeL��0ׯ���p����4E�I��Q���} _���D��::��0k��6Z��F�:{���~<�n0�Z2��uMS<�x��J�,��	ҕ%�~t�E�P�%���g�&�v�� 'Ԩc��K՗C@�9ݍ�Q Ȭ7n�Ɓm������@z���l${E>-/8�/ҍD�V�ڣF�>D��=N��&[���~^:`K�3uw�Y�z<�e1*te�i�X���nN#�S!�0܇�K3��־�D�p&���ۅ?�X�+rNq!<�����.���H~�L��|E6u l��+3"��0i�[p����qB��Ϊ�jy�V���v�~����j)cmC�m11��J+���~n�lU&��V	���+���(������[����Ys!M3�Sg�>�e�	��0�L� +8�Kii����8��[����H�F��^�.3�g_^���7
�Z�B��)�y�L(gs��{�.�%����']`���h���V\(ρ�@���.��o�9y7R��O�.'`��)]��q���M���[⯤9�$�;�䨜z]��T�䃍��I�Z�o�L��X���~zB U��O����)�y�k��(� :� +)嬭ܬ;�k�t���	U�Q�|Kz6w.0*6��L=)�~m�}��S�rQ���'J	���ة M�>�i�5
ͷ�U�E@�(���p�ջ��M�g#ϸ����N�"Zd�<�+��[�Mj��3��.�,�߰Yf{<G���F^1*g �B�<�H=�#�)�Xه5f�@��������
�@�_qY_��/�щ���ʽg-��uSnrEu,2��N��?��B�Q-q�>3rd��]�L31�'�㕪�w\� Ӥc��F�|t��>�sn dv��2-�*�4֝5�%\�I7�h�.�@g		R;�V�Ld��=�����q�x1�~����}|������Y�Y<l
�~l�w��_O��ꖤ\I��,�k#lC��3�_�7���:~ͳ�C,<��~S��Qx�����潵tElّ�%� &Q�Q��W\�@fH/2VA��snV��ϐ3�ɷD¾dI���,�a��PjR��8F h�Ӛ���k*q7�E?����*j�U�M��o�� �D>40M�,Vp]=D���i�nh,IਪQx�I�<�%��"���k�L���V���U�s+����6U�]ژ�PRh��УƋ�a��̵��K'DY:��5y�����١����C3��$�=���}�� 2�p{�5���M7���Q�][��hؗ'�S�K�$���m-��/��FUj�5���3H�jCE�������e9�Z��\��ݹ�����sn��f���m4�3�b��2��n�R�W�R��tܩ�͓.^���j�%Z5$00�V�!�C v3я�;�����P�f���3���Uc���}Q%�1���EPWu���jo��Ȑ�øN}!�ƉÁS�-�M�VA����D#�7*�����C��u
4!Ȁ��\���s�Ѳ���c���d��|�c>0
�:��y_�ZQ�UIQ�7pH�(<���]�HRY�D�֙�S.b#�.�s`I7��T�(�)_�^.ș,��|V���6��c��>7*&��\u��z��/�[6T!!)	��
��ѕ���IL��-Фp���[�b�#�AY�᫸�}��ot�QB*��.�e_�%�[O���ʆ���	�Tp6�H�才͵ޠ�����I꣼D���kC 6�&}�p	�nEz:�7��*���֎�lʑp��{{U��b_șu�]�;��e{�S��6�X^�HC���'��_��f��~G̓g�u�*�Gez7rFז�C��������
;x�����u��S�6�T*��e�;<��N_�1�448y�4g�(������;���A���a_a��1LY����S�����.;��s�Cxϥ�`_-�@2�U��9cϡ��;c4���b:����V�P�PJ��n#4���V=FXZq��*\�TU���`gM�4K��,��z�WPGmY-�{o�%��yfds2�� _ X�o3�HX�,��W"��v��n�ˉ��3 S��L�=
�w���v�gh+~�)�`�UV$I�)�hq� 4���z��-9�Yf�7�hF2m�9���_p�L�9j��?SZ�Z4�Ko��� ������2���ž5 ���I	;��4"���N�]��<!��T� $�C���Fu��v-ޠ��$�K�֠�_ѽ�]�ƥ�:��m�[����]As�)t��i���-�����G�U�0�$�1C敛���\�|Էw�*���Xz���|�GSlCA��S��C*(o$;�]l2K��;��A�N��"Mr�I��z@����s3�,9N�5����j�dщ�lxww��%S
�V��!	��ow1����Sp��&�ţ��[8d�>)4�ЖC��Xi��CF�xu���oR�w���a��2J|��S,�4�hA)A���]?��S9pm�=��}�3�����^5ېQ�%�0�'t���٘�< �jR��Pr|j*����%P�DZ�I�\��v�~{�>�ϑ������	�c�Uo�E�Y���6���m�9ɔ��e�dУL�a(
��"�;^��J5�y��=�����M�h���bC^ړ��Mŝ��!�>�s�ֻ�f�Ğ�3��>�h<(&
��c�r�׏k3����0�D(��.Q�D5��y('�MvP	��U�xmG�&��� ���L�UJ�_��d� ʣa��3����u�����v�N|��Q�uB��T���	�{�tn+s;�W�MAR�N����R��,��ig?'q$r)(���b��oUcF8r�@ԣ�AY�I���Z��v`���؎�Od�n�1�����3�vzZ(�B.�	��q��PgLQ���f-���MҠ3a�&��z�9�-�D9�h�01i/��*ܧ�}�QL������62�b"@�Z=z��p�����IpK��+��[��z��)ٻ��%s�n�5�:�w4�J��Og�"J�,^t2���{"�9�,���W2{{s��ue��Yt~���L�"��"�����[��#y,�q���\�F��yGݼ��w�{�w�po[)B�W�����뜛5��i�+�;�ǋqQm��TQ$�4��u�1s)R������.Sg�@�U;E�L���T�$3"�xA�7��(�~�j�"�x�SL��Z~�RKGrS۰���e����2*�[1�%O�y����|wN�l�K3��͸�1��?��4[�`�S��a�f�U+�ET�1(�GlF0M2����pE.c#�&sN{�S�����0biw���)32ʫS�\i��7SG²�z[��3�W.)�6��_a��#�a4�[��p��T1��]�d ?Gmԅ��N�G`�궫�d��������[9ۼF*��b}{cl\�����Z�@������O���݇h��4��¢�Pxt�,O��5�8�̢z�~cpѓ�+!�ō��BP�E.�^{:����?`i[R�����^M�p�<fa4����x7o43�z��L�U�.~[�@|%:+I��n��]��,���*,�:����V��ZxQK�u�	�0yf[��/�\��5;d*�%��߯��C% V3��qY|�@�hf�S�?��J���˰,Y�^��5�q�:�&p�9�x��6�~I@�ר*+��A�%��;�aFZf�!S�ǏU��(��/%ĬgA�pJ�B�I����ys?�^Z뉐^r�m����J��;�1���,~� "�4p:�K0� %�����5�F�t)�*O
n�vEg�YX'Hʟ����mÓ��2���B�ޞ����X��ڂ��ܛ�a�Yz%���XOL��N��J]CI���\��$q�jN�x5���U�4$q�m+u���[<��ۥ8���kߟ�X`y�.=�s�aQ/J�[_2>�㳻Oն,F��[L!������9��v�U[%�b@���?m�-+�U��Fg��śY������H��Գ�E�H�šVȺ�����Ut��5[ 
(�����[�A.�K��7eM�Ϡ]�:e�(ɶ��y��:�
��~�Z�m-y�<���^le��+X�sl-�)��a	%a~�J� ��/��]|P0���6�h�����M:�j�K�lvN�����\k���p�f.5Hݎ��U< �I^qo��S�A�Q5���[�u>�̙�i�mo�ږ"�m1ҺH���J��{Ǘ��k�A�c�u���c�E���9'�ӣSB�n�E�j�E��D�b�׈M�I�'�|\*܆C�01�8�-���3�'<E��;��?!�N K��Q�d=���OX4�/�6X�h�3����f�\�����4ǭ�Sޓ�,Ņ��w�4�d�9��O�0���)2X �O��eZ�b��C�����&3%wzVp�H���������;��h
MNn�Hn�{��_��%��$a�q:
x6t�{w*E�-�`�����s�k�����} �����@K�m�;o�߿�Oխn6t\VM��k������r9���=jA��=�]I������C��oX
4�4��7]7=�w��c���i���H�%Ě�L��*�ፀ�_��'�ճ:�.8�`^t���{)EvAl.��v�</�۳�x^[�]f��X w����쩅�4�ۤ>�Ü���/�JW�	�ڹy�H�#.s��iP4�Q��`�V��j����r4�I���բ �#���4Υ��7t|0<%6��b#⼣	x��=-�V����T���m��U�&�B(�֓�:w;㱨��_��(����$��k�RB��f{�P
S���`���Ftc�b�?A5*H�;\$>�	a�d1������Đh�����������.��}�?ߛ@�1��¼�vAl�A�������~�5��3L�O���&t�Ԭh���굠gRqJ�5�� [ʶ	�"�և�䀨UG���h��R�4>/S�#�G�r���ǥ���Z��>�Y�٥#��)}C�������iJ[���d�C�f�*��Ux0���ռ.�o�O|v��1u{UH$�p���T��68@#�?\�5@����o��m�0��J0�5���v�8v�h��/|�±�LZV	e}�׹�Q�\�{@/��J�L\#�n-t�^r���m��N`9��}y���k�O�mh��F�Ӈ�lgL��#Q��wn'�0���6����X��-H+���� ӽC�c-��/U�>�ߘ9�6"�CS����{��É�~�~��]��$���գ�HxMy�1�79��w9ZL��wF��v A�`���QA����Qf���n�)�RF�8r.�e\z?�f�;1��Vjn�T��t�4��)�k��{�����]���t�l�x���L^���D%�#H����Z֔�sNPx�����,[=/ �h,�B�F������p��,�70�%���g����Z�-�v��,�0��y� a~�?��������4�T�`٫A�=��t��n⚪溥���h+g�`׉ab��,o�	���묯�@=D� &C+#�kUW,P�Tl�<�뱒Ac,����w�ڟ=8A]�!��>�H��)�cm�

����197]������{xǬM.G�&�}/a����;]0��-�НJ��op�әc&{��	��`�YM�#��v6Y�_��zsYg�����&@A�5�w@:<�e���l\|���JrlX�<�1�n@X��Bv�&�7j��eK��B�̧wA�B���� ��fZA�����5���?�0�~��޳T�R{d�jn�3�����'M�u!�{�,{�%>��qx-p�x/��*���k�Vut�~�Ҋ4S�2\��XKρu�����e�OX�J�����HM���~���9�p"���䴪+=
�E]{�}f�#a�Ld�k�
f�Cy��{$M|���X��]g�fD��o_�KR� ����h&���)���+�#�P.$ցr�yV����eٵ$��K��C��|X�%v�u(�y�������r�WS� ����A�AU3�	ۣ�>���,��[G��,]+�h��V�J�̰f�i���������)�T�t�\F�6������X���ջFt�Pyqu��Ӎ4wA���[#!eY:���M��79iy���&��T�[}Oom�@�Fb���Ƌ�,ҩ��^���q(�&P󥣒�{�!�1��w�`���2gD�$�%�}��su��զ��6� XA'��d@����߫i��	�8R�m[!�6�3o9#[q�G��w�}ޮeL���ׇ��Z���ˡ��O�y��17�\�W��{����K��ok��t5��П�*����c�����8�.�	�����Z+U��(�8���$�񄏃G��ٴ͐�"�n�����U�?d�V��?�<��"@���9�a.�T�Y6`��Z$���p~[�7{�*���Ι@�C�e9��~�P�ϩ�BR���f;40?�0���ko�UL̏@r�'�Y*��;�B�������-��o�n�x�]�[%.=�|�}ou�sX4��N�2s��c���8)�����������Jy�R37�R8��LձUE�Q)js|�-��i��Z�o��.2)����1N�=߳[�#�O�3R}���)AJ-�1u��fj�4E���{�r������Kl�:M�N4A�j�N�a�ב�&�� z�m��*WW�	_Z�$9]e�B�N�Zp�̐rO�V+G ^�>��"y�+��p�w���	a���&�V����\0��jWZ��ig��G;/�i	�@��d���V���ȕmP����vY�o���)%ֽ6c��q�g��!�"U�K-A�F6�}G�9E��{>�������(��s�eݕ@��b�=�i7R������ΧT�}�r�@��"���1}�/�@{j�i��
��]|�n�		�ÌS�kes��gg˳E��3���>�a���ţ����k=\��Z���Pi\�Y^Yb�,��5Z�}�% �	|�[4tm���̃�IGH^�ߗ/y1�]Tca@Axh!�Ɗ���́�����I���'X�rf^��z�3l���JhN�:��'	ߌ�:è0*�ECa0��(�Ā%Vw�t���	x
ź�C8��g Ǝ�a��[�ۣ
i���7nhe��R�;{�@��3G������(49utw�#d0�"�C @�����$�C|Q�r�admlpr��w���&�n�r+[=ݭѷ{�9҄��ȕɉ\�L�e"^���r��2S�F.�|sKKǭ_,p�))�R�C4������s"��Y')� i;�6#�i���a�)3�0��O)�'��ly璸��&]+�$�H��_�B�i�����
l�
�x�����\&�sCƢ-�#��G��|q�r"�T:���Iư��8��UW��s�㷾���&���NLr��֢�TZ�� ,c�&�Bf�+������/�>�`)�GM������I-�O��U�
q��d7L�����<|���4��l��E�2�72V����۲^b�fvT����� =&v�Q|�V�*����Ĥ�8�m���/�גX˧x�:`�
��/*,!�Yzw:�t`V$٣.���ؕ*�&Jc�mft�ʗTNn<�!�*��Q?괉��	�������
�V�	�0��;|�!ݻ�O���T͒[���/��9����¢=�y
T�Z����G!�i&����ǐ���Y��<��۽�$�9{����"ʼZq�#��޲�n�=��_�����]�&�䨙Nî�_aL���x�P�����#�).=��_�>'�7`z�}�8��ƹov)���;���*{%��f��^EM�����)Ҿ8�|�j�[ߵz������
M�j!X�[E��r��+(Z�݌�L0��J7��1>�sa�U�~A��J%M��,9/�����~K�c
3_%�d@fP$"G)G��!�g8��goMt��k4;Rs4�kB�w~\�1�	J���������l��-�-u Z��%��)��-�����jH��#1�pP��2�~��A�w��8eXG,\��$w+S���0썃><�͗ꝋ[j��B��f��f2mE��!B�X,M8uư;̋e�o��2p���;�i8��0�7?pN ���6�.ۉ���%�ٯ���i��>� -,�����wZ�����
7�M���Kʵ�\`�|N��C��8�"a�İ�=}w^$��������wW������$-��X���J�PZs���f�D�����F9�6-��C�6�vF�[<먜��8Xtoe�~�ꍾ1�ɮ��AE��W۪�cSB/��_m�0���}�7������i����X��2T3�|77ImwG���ƙv]��jP��%pVbɳ�c�w����
��n�5�ҩ����]ɛ�F�<
:��+���L��$��J3Ϸ����}�OQ��5?O�g;��즔�D��:!]@��Kzi]�v��y�)4�ͽ���yO9[A2֫��g�t�2ؿ���@9��b~�Lʀ�+�\�`軮��)\��E5�JMό�����r��E��Ea!�ϤK��@��L�Ӆ��wi,V��$����7Z�N���_�W2��7"����6<*����Y<Vޕ���f�1�/�[捖[jOu>JÕr���{��ִ�J|U H���,��/�1a4�-�S��>��3m�o!Ό)t�������=�UGv����#�QPB���W�	��Kl�髮�z����6���~ӗ��5`���� �/�u��@�Uɿ���g$���R�#�.�$9�?2m��P��v6���֦��W�oDJC�q�Oz�����s�w)|�53��\��̛�GND�-��L��e��Cv�E+�"KLƾ:�K5���fjר\ZM��=`h-�qҮ��,
\5i�D�1����O�C�̄龩��:}�h�y���"p�m��r��������uW�)�@�q`5!w���ܣ�}Awǵh�xSj�f��[��k�yH<���1���ī��{�&]��A'w��
�v�������M�;�^T�v�;�d�>�͸���������_�׎��b	k&��P�_6�_�X.R�Z0RwOwj4r�{>�D�1_P�����3���,MS���i< ][�a�1SJ�Qh��~J?[g�t/7�H�aVV�5Sw<�yQWXc�̓L�72�*�������M�5����qg:�/g��)f:՗��R�Yw��7�sp�*��J�#� yR��u<�P�mTuW�S	!� ��==���-HO݈uqNr*O�����h���)\��ԽF�my9��D���#��j�퍔D&Ó��9���
K8�����/J�����W��T��S @G�^��_��c�>s��0�!8�,2&�Lˊ�
��[�����G��������"����.�����FL�*��y����S��h�ҳ�-�n�o�7�k���&�=9��>�K�~�*`����$fJ����D�/X	�D3�i��]ܺb(JMJ�b�^傘nd�n�.XV��SlIM�h0YWNWKbG�8F���W3:N�Z+������2�5m�y���J���&C�f�ç��hL!�M4��ٻ�0���8�T��� ;�D��͠5�E��)`,�0�o�Fi�o�oE�W��|,�<B�i���=;�A�.�D��Y-��c99O$6�?`3���yg��4�%�lZ�mul�ԝ�^]��t����(o�!��p�3�-�H�c���h|Rs�.Y��yΗ?�h�W�B\,���
f�+54�w4���NM�՚.78��j����0���j����tnU`�'���+�+$���z1k{���8�0@&D�ҚA�t�[�r��*����
��5����ٌ�S�����tԓoS[-s`Ic4mO���3$Ü)2���bk��S3E0Q��9I�$�&f��l׹K����{!h��~Qe����w[bJ�gT,��c��L��"�fq���������l$ ���>><d��	7ʳ,cQϰ������T�� � � 	�2oo�v��FXs-zf���%�`�=e>q�$5����;�&rA퐍�����[7�����C���A۽~ț�c�00����+��I���?
����?M�^v&��Hn��g(�4���Or�	�
Sxv�߫��}�\��>�c*���Xn@����N�g�pI�oP�����W��?���4��E䶐h-ѹG��C� ሺ�AI$qr�� �d�c�'Կ�V������aӲ����%5~���#j�
L��Eh"�~nUl��-�j�<&���a�e&d��+�jQ�D7��U�Bߟ��}��z�S���	��2�ic�:�%A���2xU����>��P�FC
�������y��W%u	�m$Mi/��{��s�wy'�fMr,�^M��yP�TC�!/$����/g��t(ʙlK���~:F�˲C�9ا�o2I7�+J�i��{	f�|� �QMQjD��D�ϳ)^�ڹ#�%\��)�u2��x��K�}G�E��a�6&�gͤ����Y���؋1���6�ql+Zp�q��Ns8w����P;Hav�R/���G.�ձ- ��C9�ɲ���1��ڮ^�Z9S�$��])��? 	�yS������ ��R��L;�(R_m,�{a��'�EM�]��	L"���z4���/�k���]˝F�m��6� '�ɋ?ʝ���L0�s$e>o�h�	c�*%q�'���]a�9kK$�:��2l1����z-�(v���J(\��.�~��c�W���:�2�R�7R���E��Ʌ ��hM�A'�tj�����7���:	n$���WS��b�	�4E��}��]S�`J$5W.8H�۫0���PP!�V>I���K,-B_�Xboק�c�wa S�ټ��X\.�Ml���~�S*�$��~�}rX͎{�؉�4.��T? �Z���3f�=u0�}����\jEw���g獐�1�Ue���4Sm���T�s����`ؠ
�W���Q�K�wc�=j����)��J��4\�������w�]7p:�m�Y���Xѩ�F\�{"�2��e8��t_��?P-?�ls,!+���V� �Sb{>�6�#��*�R�<����rܬ׵�D�VE-˴��Z��=��"l*ix�^9��Q�fG�<1���ř�w��>��M ���,N"+�Ӵ3rJ#���k�!� �6�1�g�'���Iw�2f-�˫[�-SG�~����*��1�PI#�ī-��H��V��0p�+E���,�,��Kr�_bz��`���y!K��3P�;�Ca8k����c�K���Z]l�,���M�?�/�!����v�H�䌋��g�<8k�8r���C\�]��a��k������:�B!�����2��*P\)g�\��C���l}���2�LG�Ĕ��9_�{v��:�`���8��%�|M��#��۲�47Zɻ��|K����Z^�n�%�ec�឵�7�,�8ۺ�����/8�++!�q�c�eh����%�!�RR��|J�h� o�����@�60*���k��pyd�"���3�ۭ+��i�]Z�2�DTu��a����5�굋��W����~Ym���`�����`������V��]�L�ó�k� �������fw��-���[w��������^>�Z��4�xe��%(=�/n�P�dB��%�F�\}�~�m��(���̚�.Ia�!$�ʒh22(t	�C�e��D�"K�,�%V�ڛ!�C���g�owGl`~�
�+�8&]���� R�߂�/�֭�ݹ6�:����!}��䧖3�٫�]��ޣz_���`Z�-0�loE�)���\z����:�n�rib���<���u@�O��V�m���!1u���uǲ"LH����@f�_�]�`�6']-5����`�N�_֘Q��_N�Ak�zkL\������ ��W":>��_��s�6z��Ib���BT������LK�x��?ܮ��'�#�ZG2
��ϔ��>�Yw��t��1r<L-R�l
�J�ZFdk�kYE�Vt6$�俤�P:�;��g]j���]X�b��1��Ν�-��*\�+G�����nΖ���Y7�����;W�A��A�w�����.��io�-X�)Ԟ�o�цƣ_.8βIo3&��n�˯�$^��,����?���D����]U7��~��ɠUR�\K��u=	`�uұ��N�������C��{�6��L�ֈWn���-�Fe�Yh5��/P�����*�Э˝I�Y�.y�6�u�IM�\��,�^9?�4��x+7B�|Dl��.S7�oSS�j�o���%!'�5='�i�7v0s�a���4������ܯ2���P��qF1t�RDN�(4 ��}&�j0���=	q�1^�ԇ��׮1�Fa��sɟ1t�����ܫI1~��s���Y���٧A�l��X32ڢ
�QӠuT�o�����% e�^�1Q�l)�u��W�F�(d�o���O�t�zӫ���)��j�PL��Z�]���������T�����@@(�jVmRJ�O�v�ӆ��'��Y�nH�wj����~:��h���e�0���_]���v6k}�q�
�i�@H�P����� �8'?4���s�h�)��i���Xj#w�z���|���g�(Fa~��(Vw<"�d
��-�
����LPb��@+���Y������1�3[���_�\����� Y5<�A�B�ϬE�g������	m8�1
 �JB^O��dU^�;n��r�)@CD&a|4m!������U3G�B׆���g�t�%bC)7l[a��y5�x��}�x/���ʏ�d"mS0��U�� 3�� � A(��Oie�
��$�Lf��e���gj��y�&:B��r�9АN-/�r� �cO�rI�U���]O��|��U\c�gS��Ŧ/�!7l'�Z�V|�;|�&��L ecL��/��>������|�\2�|�>^�Q�R7͍���J�1e��h�(�H+a����>�����dN�jr�Wx�tS�u"_�w�Â����#Ta������FI؀���]�1i6W���O�5ɬ����g�4��c�N�	��^Z�.f\��Ҵ��Pc�M�jq�0�yw\�_�.l<�AV��#�!��#{��i��f�:��E1~Hv)�������P>Bz{F�&&�#"D��'�u(����#�elT�b!�	�R�f�.J���L�ff��q4����Ǫ�]^��_����7�,%�FI����X�f�1w� A;)"ui����k<S�Է��S�U}3�������ԭ���e��쮝���ؑ�!-�<jB�c��"�!�bE�l-��8!�w����I�s���f�Tq��D�=����@�ª�� �
avΤ��Q�۩��VQ�g���z�=�M�aAK6�)NZ;Cq���K�[Gc��Z��-���C�Pƥ��(;[��-�R.%XC!f�)2{ԯϣE�� Hd�`���\�$��'��FFʽ�A�f8~��<����� jŻ��滥�v< �ح1�)��L�������B���<|q�̤��A=�W��J)�U��u����� �ӣ��A�n�Wv�|�yT*��pZ�N�͆�T�<�xR6d��n`����V*Я+S:c�޸ؙ y��%�� .���g�k���0�$����P���/|�8�V�9�W�v��&�A��6�/���e�����o%�/Y[�ʤ�l��Ͽ��4�@������d��!��T=�SR�g[A�g"
�ޱ���/m�g8"�r���A}_%kY���N�0��P��<�=O������������A*����G*|'+Y�7����Y��t�3�x��B��w�V ׍+V�Ӏ�U��F��k:|�A%nē=	������w���ۄԗ*�9�v*ـ~K���}�<�9��մ���jZap����������Qlïs����/8ll�&�}�I�M���CȨ��"9�fM�[ԣ����6k��#�2o�H�θE<�;b��C/+��clQ�з�G'���"x���t�&E S��ߋ�[I���U���R�I������^�)c�>L	)3Ay�aY�nQ�������RM��7�X����Z+G�n�7�!^U>9�����kcf��>'�:\�q%u���"�fOԴ�\:�=�LWz�8-�ɼÆ�)Q֪P��bd�n�n�x���*н��B ��u�#	 �-,��"�EV�d ��O+e>z䭾���.��j^D63�M��J'��۵���.�t�s�:����{�>�Kr�=���/��g���Ո@Ҷ�3������p^<�E�XmT�����󎻲��C����?�yHwQ~�fC{6��⑉U��*��� ��<������l�.���*�u\?E*
��]h�b�P3���{F;^�`=�9K�Q���h	�5��y�a��^̖3'e!$*�'@xշ��H�����*=�j�{�^+q�*q!�mqDw�ԋ�7R/��lӰHa���/:�\H��� ���ٻL້�^eFh���'~����{6���C��G-Q=�I,�st�p�6������i��ɾ�������)X"�5<��sk�LbO_;�C�ĆGK<��L�Τ�k+j�e󠴬�='�����tva�d�ѐ��whA.��UQܒ����05k�W�+��_�9C�:�}���(w{W���p�cX���9$���bq�ɡ�э�a5~|�ʾO���~P��x&��j��V�	N�j3h�����`bZ�w���O����2�n��^G�f���,�ʜO�膺��~u=Ƣh��BD�9x	�9.�^��~�:'���<f�4jcm
�T��~f!��[l��5nH�2�"�จa�[�"��\��x���o�X�~@��,�v�i^��At���	��#�����U=R�n.�����`�{��3��fX؄m�+�����8�c���s$�.��X������u�IJ�������Q���6����j*�����lU�ӄ�C(�*|B�KM�N?D�����qr��)+�J���j�a�b"`��I�tK!^���:?$�h��$`�� ���|ah���{��$��g	�9?O.�
����_w��Q{Y�{�Ɓ~��ڪmm#2�G|��H��P�v�%iL�K���F[�P�Y��se��'�Je~�T�+AU�.��(/����w�EK�J�V�vM��S�(�g'�a|�
�-h��LV���dY�zy����{�ɤt��M�9q��@���
�ۻO�l� �=UφR��!TŽ�
�Qj��P(F�t�TƼ��M>}5+T��mS�ߤ��� �FM����,�RK����/��������Zf�߻ڷ_ ��fh�PE�h��Z��,��Q@����R�@�<I�͏a�]@�23~+6w2S,�p��/���)OW׾,��V�L�)[��QU 7D��XU�u8[��0�T�Z�rZ����" ,�B(
s�lꃁh@�ell�^ �<�qs���T~ ���"bnh��� ���}Oƨ��@�K8�?�7$�~� ��1j�m����M�3l�I�L�y+߰�˗����z�\�D����[D�s�1��=�Tp(�q��"}�}%;�#��8�����0���W���;�\P��KF��N�.����p^T?���R��}V����"��qd\{�0��B��G��.F���-/G�_��5X�ظ�O����K�n��Rq��e�?��3��#0<c�����AV����q��~]'����/|&���y���'Vm_���������|��ۇ!�ʔif�~�ivL�����( K(1�J#{%ߠ�j|3���J
�Q7� ih�q�3�b��wK������V���o��m��`��m��ɢ��
&�
�<���(D=S���1�#�>��P� ���2�X	�˼��0��b/|cC3p���wͪ|�kXX�ϐ��!�?�L�������X}��8	d]p7"f�]f{f�S��+{T���ܝK�!(�L�	�z^�4 ����������˷�i�(4B�I-,9v�:��>"Jqȟ�P�V3�%>zg\��az��S���q��,s@8�~����cs��(�m�Ij#^	��z�D�꣆�����Y]���~cz�^I�B|۰F��)����*'��0�b�(�q��lU'���$9�^#�#�Ã�=sq/�Е����V�>..�dU7-�lɯU/���o(����4Q�YW(\O�]�۬�䑆*E�3\��Ȉ wc7`���N��/w5G|@��օ�.~������N�~���*E@�$T�謀�F`�z���Ie@-aWO�e`|(kXJ��tr�;��W�5G���2��<�\����t��m/y�ЂA?�ZMXI s��1g��_Yz?KN��EDj��<<0)��3Z+E���뤖~�I��r�'�o��ʋ�$���8U�bG�3��Od��p'�vaP��(ߔ�wtݗh��9���)�o�Z�� �A�p=ج�,��i����lx����렛�`\�h S�N\E�0��7�ڡۦE�r}�%K,-Q��Z5��6c�@�;��9ңq�k�,a>����7�)���傌�]�7O+*���L���sj4����])�ސf���lVꗋ��������v~Ź=�tg�dQ�V��������t*�n�)S��ަaא��\��Q�Ŕ�����Q�D���y��#/L���nn��Rd��s����U4�@��_
���w���,���G��(�#�����Tz�=�N�[�������Q�-�_������F����YV�5+�{�������!�M�����6=IL����s쨀`�Ԑ�#�ҍ���RE�.|�Ŕ�������QT�cS�c��8qy���5��.��o�Evq�}��@��H����s���t��]P+5�e`-����|��U�Y�֐��l|�R�;c�dR�%�n����i�����/G�(�h�b�r��bDPFZwB�xd�.��x;�y%��.I�Ky\⧘�w�fy����-�Oq����� U��Ef?	��Wn�e��֪�#�xR"AƲ,��'V�]���rL�sU�O����ׅ
_�{�k�v�ބ����p.|\4l�j��D��hCL��s�Auz�����b��S�t$#��χ���J��
NXq�Ү
VZ|7hE(���ʟ���8�l5���� ��/���y�c��޿���oМ�<zY"�v��INO��^��e)Z��*�9�̥d�y��I1_lW�^a��ص� ����~��!}�� u
��%܅>�?���*��o��@��\`�/3�qr���Ԅ��p�_�V0���
����x�o3�?��΅��:Ž>�����X�[DT��2�q �H�K�	iytA�ϛ������B�B��ʏ��L�QQG�U�Z�&9�[U��{��hŒ�߼�Y�H�t-�x�ѱ����s���_�����L�~˱J�J���_J�w`K�K\P��K�ԡ�2�Z^��&�����4�w'�D@0;�4-���S���c�����BT8<����g��2Rz��{�X�_�hᾃ��ҏ���S~���CF[T2��-�64o�Z�v*��< �$J߂����L��8bzI)��� ��Q�$�����w����u���Y	�e`������� �KY��__�R�B�?.��mw����j�0�;(h ������]��_m�wko ������}�+F�-Һ䆢H����e�'��<S�g��{�c��D����J�v��՗0����V�MG���"��1��f�SN`�-���n�gy��1���&4z$��5Ęv��_�sO[�� �#x��0��� w�+�܏���d=iY�51����o���O�>XY�}G�1��y��+�]C�V谖̴=�$9Tt�zb���S8C=�@'��_\BI�X�X����E��-���تł'���b��-�Z>�ϔ��������P�����l�"wI��^�0ԁ��dC��ᆯ����� Uߎ�n�~���ߪnܵ62���c�b!��?)P�t6Y���N��p�����Ls� Mӗ��@(u�*�;�R� <:[ 4]l�����Q&U� u���|�;`���}AG����5�I7�0gȥ�u��K�l��r���U�[�d���9	�CYg7�׵��ݛ������@o�Ĭ���m�zY�Xk!bDN�>ldo�ϣ7h#R���u�N�F��z�<i�[���u�!�Ъ�W}r��0Q�u��:��9՘Y���W̨O7?��'{Z�˰v���W{y�Z;�Ȥm��D�Kx��{�8��	��LtE���$V/��
<Y�[.?�GrO/������x�$���Y����4�k�|��	W��K�ɑв��i\�U�@c#�����R��c�~��T�Z���(`�����8�V(�������:$[���g���g����QO�t���0�%������2�th� gE4<N\P$��k�/,��0&F.d'i�?�A��$��Aq~����]�1?6�h]�v���,&�ڵ~c>�Y�U%�Yq����m{�r�z��:�4�{#Lhv:&������@i|�m3��,�3Q����tot���m�t��k!�`���~P�����L�I3KRc�d`�m�	�[@.�*LB�"
��M��l�g0�O�jb�>޵��*�m�	|꙯m�#r�5����~&�в�dB�8Wc�����g��q�9s	����������F��Չj[L��.���ZY�OZ�����m�@��>��K��s�`!RU1����J����q2�����z?Z�#Uyg��G� N�ɣ?�n�E���F�U#(�mLk�ܚә*�"�H���a\΋Q���K"�	�6�V�DT��g��	�Vж�i�%[��s�������j����­�t��CF8��b��$8|#/�����a�眒�޲��.1��O}Q�l����+�%����6��®t�_��V'���"kHu�(�[�>?�%��n+�q���,e��3D;И��8��ax}�p\Ǆ���=e�eT�(;�����X
���4��LH��v�� _��)��1��Fx+H�1��W���?�	v��?Ay �Q�As�G4J�G��P{��A����B�#j�u��1�� �t���W}��4�K�Fn��i��4Q,#�0HM����(�������wg��	�C��T0Oh!e�~����X�y�l[^]FV�<`��u��)x�(}#=֢Z���Nq��2��Nqf��� ��_����|�es�蹦�CkC3��&��f�8G�x��M��8�Jo�Rvd��5=���U)Z{�UH�|�q+��kg����^�36n�gB:c��-�r�d��)�{�Ѿć�$$�����L��a�P)�/����7�@B��k\ڽ�����g)6Ɉф�7���Sr'yJ��,�.L	9&�J5z�ܶ���6��%�4�=)��T_�M��@"����ch���,P2��3�ދ<ԅS��0�,"\�S���fjї�.��������d^�/>����{�z�c(��g���"#QǨ���e�/�h�B5ӗ��ˤL�C?
��e����X�f
���u(B��H�D�S��X&��upi��*'֕�[���[�5^DNB��+��U�
8��鐊yבP��<K ��#I�ΡF�&{��ˉ�[�lrrD���#���R{Pݒx�Id{;��t��ud(H��_��g_'ld��ynl;_^��uj��<��	)�l��� !T�#� �C��b�����Xï"@�F�S��p�/��"���i�� �|I��	��.	��4p��:���_p��f2/[���SR���>Q������{���ʰ��p4�8��^�/�(=��v�����P\.��%r$7J��A���-�IR�(�_1q8J�~����Cq�4����jg��g�9��^($7*�m��BG-b��@��.�_g��$�t�j��i��w��%���Z\��,��A�6��~�B�'��f0�X
	u�S-�*
M6�B]И}�w++1ܼ�G�@�]!gr�A���H���X��TWivU%H��%ǡp�қ+���F͆*v~ml�x"v_�!��[� 3��+.n�(I��0��%.��iP��?s�0��۪?}!ϯ`��`���z��?'C����꧓?Q�-=X��Z�p�j}K���R9�	�����?���Y�BoS������l�"���gh���h����X�u�i���@�4t�J�
^l+BM�&��R푲 骍�N��z��'�ŝ�|G��j�+=�2��b��c?VE/M]K�u��>���vS��/4�o�5&R��7�e\������	�W:�+*��8=�	�s�x��%����"�8�Ͱ�k:��fb7C�	Y���%�.�xnZ���^�5�G
��-�*M��.�r�-�vU���0�"8��+@���n��g#��@��n����*�����B9�q�cd�p#��W��c���j��!������Ƃ��8r�m�_�b��(q������g�*�x;V��!׏=�٠"i��rp��E`Zo]=���~/v|p��7d"��:�����Bx\��,��6�}��Ϻn�ȭ�i�t|SY��A_x�#�A�Ɛ��E,#r��qȱ��Ez���(-%�j���8r{����Ĥ�kԄW�l�*�U�P�G{[S	#�Q\%q�#�(^�kFA��t[����>OS�}��A�J b�̐K��(헫�x�h
���UQ4L<���c��c�&�;FF)�@4��г0�t"����s��8^CY�oy�x,�s����m���>�ZD�\�(S!��2��;�i!H�LWe�	>��k��F}�~YCXs���둞	��}�2�\��?��CԟL|�7#��-s���&�EZ9ۮ���Fv�	�(���Pw뚰X@���)�^�!�MAUL��Rd���}���oF%��CU�30�)����}c
�i+�E�)�t	dI��\r���mr�a��TF�f�q|U@�R��u$T�F��Fi_��ZX$��{r�h�U����_dj�+=��V��_2�⻞�s;��W�A�z?���i�l����a���o�0;�����"v��V� 4
��������#~ϗ�l�Y=Ѩ4���=�)F:7�u�g�<��f�?��X����$��%�r]ͫ����m}��W�DŃ�<s��(�OMVTa|� d�DXi�N�񛪌��g���s�f�!�Ôf���pJ�U�~S���HTc5�V��^Y$|� =ɧS:,�9顩b���Pu����_&���ɝ�q��ګQid�LZ0��x�_�8$3͈n:+n�8}�>N���Tn
��$`+G�	���:�Ĥ(oh�R��7�_)�R�Q�l�3$���M4i�	�lV_|j��-0y���jv�p�e�I]K���R�H�ٓ_�w5&�q"B�8������Z-�xl���tVOo�DNv;z���K[�B�=z~y<�ʌ&d�������������ܮu��@<���&ܕ�m��A<�ѿ.n>�&aG��ߌ����?u���HQ,e�,>]�����:7�j�E򘀓�Xdi�����{���7��J�M."�}Ưш	���#�E-��Q����C�b
d�'��LB�a���S��N\)����Â���%�| @�N �XMB֙�o��}����S>�Ma�v��K������Y�ÜTWe��WO�S��T�ɝ�㡒��vIG�G'FQ�kJ���R$?Dj\�b��S���i(�#F|�n��_����NqP�N[�ȓ;MjKB��v���\�ԣ��NҰ"{>�|�e���+��NC�OKC���mRx3��&��h:U}wta��l}�<�T]���>m<Λ���r���T̀��)�{�-i�`^�ɑg!��i�].aX�*����<�_���H�J��/A^�(���|l�:>��(]���,5omt}	n�Ur���{�ڠK	��-�|�1.��b����?j���R/}L����S��S�Ϯ�}}2���˕�����:��U"��hy(��}*�ܟf��,b�� d(�?V�@@Hlxj���½��/�xp�J'�{P���(��e�\C���|"�SF2�XMGZ�<H`H_P�H���ڼ�)�~0�8}6]����3��7<&,��C�sB�f8O��-���_,��W<��*�b����p>��'>;p�Qr��JP�s�vx�NFD%��_NzҺ��2�� ������� �Xu�"6VT������,L��u]�E	�A4���ܖ5v	��)���l�gkȌ����h��%��B!W�v�M�#���)��������m�碆6r}�Pą<�)ړ�=��c�@8�W����j��n>�&L���)xr�`NJ��iD?��B�+�ޗy%-��u�k2����WG%ٻ��Ţ@^�'�pB�K��a�g݇s�K����Ί���^b�@tѝ��U������˫U,�з��6t��z��	a�����Q�(I��d�ܺ�
������h�S�����������򨰰��׺4h�}V��Lע:>�T�������d����h���D"���G�Q]�t�g�v���Yv�C��f^�x9[uKW�GZ �����g�s�Q�J���}�",��y�T$%8�Dm�P.��i��0aBo����?�N{]}Ӣ�&�_+���.'�p�n������ۢW!o��9_Dk�F�|A'�(��v���_����Ko���֦4�,�����ˉew�$<�*�_��3\��^��S� ���5��i301	���&�/Aݞ�rb�,�"��?cB�ގC�%U�bE`�C}�	�v�H���4�0�o�$��q[Űo��W�3��M�" b�Y3D���F�H���[OU7y�*(~x�z�Pb 	2}����I���OO'v��m��[j��� ��]���I:��O��M�
1�\$��Y�\�2��%�µr��L$�Y�Tȗ��j���ZN='��h�����]��2����A@�脂&�,�7�°b��������N�Hኻ�*G��z�g��x�Aj��.���z�����ju���ڍ.Q��5#P]�P7�>�=��b���(y1��v�V�^�/�����Ɔ,�f_V�	���Z�@B�I��W����I9.�XR��(�Z�~AD�x�{��D�\?N��k4�|�a�� �n{��P$��7)�ߵ#�����-lɢ��!��UX��CA��m��X܌�ӆ�Fk+������ `z��Iw7��a��[�Q�qa_�Ŗ�D��D��ђ*�����o���~U,�f	y��I��t3ջ!g��1�Z@��(r!����b������l��k'Ԙ�#�{�C]�&ЈY�4p�̝���K UǈÓ_$m�����d�e�*��z]ާ@���e��F8�UH
TG?�	��-�7b�:Er�f����Z��7nb���5���L�D�LK:,y~E�l��M&N\�4��wh`8D�A�D����<m�InE^ԟ�_����$��m��{x�1����8��e��q҆SSl����>8��3�(w2�����c$M�EO��5Sk!��=|���?��aO�e]�K�0����G][������Y����KcSw�(CCG~�J,q�Á7�Z�\%�Q8
�m@���@��e�f������`���e76��nj��خ������E�l�{@��,�b\O���?���?� �{���P��gV�e�\�%�|�m����V�֥�.Q�DK<�P3��%'~Ώ�GS�ʾ�%ޒ�����k�� :8̍)��K��sl��z�����X<�+Ⱦ7y���lhX���$�)�Eq�-�P�����Bt<F��!(�p
�N�V��x�8'=���pm���%	�x������
�D�T�.���Qʲ��3}(b��;�xN�b��ZK��3Q]X�R�}�@JK0�򫯡�F�s!��6c�9��O����q����1iU��M����vaY�5A�8����V'Oh'=E�)��l�LJvTK��+���G�P/e��|H��2�
w�Ą���"S��9/z�x��7����W�¹L� (��?�z�R�R߰�*���O�8�6��D*,�١��A�uhl��}r�;��n3SQ��Xӻӌ�x��j�L��^�NѺ�"�=7����ꯏ�M�ޡn�Mm�8�EńW%+��2�Go����D*�]�k��zZ���2�\���?����6�+e����X��+x:�����؀
wvs�A�m7���b���� �)V��^��Ւ�UL/@�]��J	jz�B�\�޸�:���#�������D��)�E�<�S�^�)G\`�~�������'���-���ӏ�j�.���H������((<�9�@�>��8���@2�󋹒��<�`"�	��|���������6%�pL�J[�M�+�Dy#���3y���]
 ᢁ�6�tb��`���Yh̫�cᆠ�JӁ)�jF�$Ж"Wy:�%oh�h�Ԟ.O?��m��j1�.��bY��iC1��[.v�j�DF�9�O�eE;\���@��M[-(ſ�t���i��]+Խ6�r�Ns��a�ʻ6X�|�EQ:",���s/��JY�����gbc�r���ݶ'���a{��x�b���p�7����f��\�����{�w�4�a����<���y��H	�����խw���?�va����ǀށ؆�x���9�7�³A���5)8~4����\,��qƆ�1�a6����
�d1������2��~�Ɩ��M��'��rG֜ZH�,�U�8�(�r���2�!��m��hk��^�+��E�N
軕�������A�i�,�J��n�e�ə��A�®O�"V��|Y���e�>s�A���;��CN�M�c��a��Bmhet-�+"�������|b�o�_෋ut��i(�nV$c�64�`1V�6�����wIA��:e�$]Z�J�#i�Z�1��*e]�m�^Mo5��ȗ���W@�,h�,���	��3g��M��f���8��.����:�Ch�\�l��z��f��0�QM�!��9`I�`����H 0��_?c�����Z�������F4��dCHg�zg�֒8����$���| F	�V���ߺ���Dc���{�L��� .s����g�a��ϊJ��Mכ&G�˭��13����f��W���N��`���Q����4fb�6�3��ź�Ds�uhˉ�"_�_�����k�=Yru�K]c���G�U�RYq|=Jt�&`�d�YN��c҅?Q<'�Ì�������#?�� �| *ngMN��d��c��((�l��m�_��ǔ��Ų
�#��۸�{�H�d�c��	�!������մN�1����%=�1)���[I�)@5r8�m��i�84F��8ʏx��-����9>�����L0���D]Τ���fRKa#E2���Q��e1�[��r�d�Zi�u��͜���yV�����U�Ii���B����И��4�wlryzm�qe�^{�����0ԍelħo�Ř�GLyw�,[��"S�|T	��j�Hp��D�E�?�-KO�5O�q�1�rU���h��=i��[@�̑�)	�����<�a˛� I��m`�i����p��Բq=���%,�+�JHH�lπw!z��(��?�9��PG��y�_�N�גS�򉁎�3 n�Z�����ԷP�]�� �^�!��fb8��m'��ls��Z�8J)�&�h1gpi)^w0_a���3ll��]Ʌ��	��_��K�N_�(��\���`�b�*�i�Y򚖽���Dް�f�)c��/�Ơ���r������!��p^�%�;�-��Z"`��ۗNU����.5�^�5h�N�cV�Mw��_�A��Mp���~B�%o`m�Hk=n�%���rK�m�Ɯ����uz����n�j�	���e��"����{�4�(�$�]���&Ot�P���_(p���&�j��gB�QANhjIF>Di���~��o�~`Tig�Ň��d�!��\tKA�B1��j�E^O���������Z�^*��&���?Okf��lF�&��³B�M��#E){{�K�Ļ�4R+HM�
�d7��"H�t�I��hP�9(K�!�z(��b�O'@���d��ƶ�q�ja[��Sv��vѠ>���$k�}-e� ��Zh5���WP���B+M�Drʪ4=@f�����i�o.�З��R#E\��T�Hn��:ԙ}n��"������q�O,1�\$�s�X�E��D���j��<��7�}�o^�7~��Kt�o8�c�2el���C ^���f�^ᆫ�<k<঵��;�NZ.@�˭�k�gB���U��[IIq��Y%��7��ǥ#	_����}�*L�	��ܕRQ�{�������cmͯ�� �z���]��̫ ��$+o� ����X��UAM\�ܿ�68x2�hZ��G]�U��]נ��h~����EG}�G�p������� |��( f�_U��A�1�_jC��|�h����%U��B1�E3OrII�@��̸,ol��G<��M�"�éN���4<���O�X;��/\�����,΍�]�QW������]h��:�gz�]��U?X�тP4U�-uo�]�b����z)�.�_���� �p,�2I�4���۷ѹkUt�>�(>F¡V��`ۂwy��v��]�l�pC�{cA�ʡ��F�e1��?\I�N�����}4�w�����X$�����9��dU��[\ፁ��Ȗ��HCL#�+� 
�,�"[��z�]l�=;��ir�X��d�����m�҄xZ�����O����5̲ϖe��8(2K~��\�{��s�J�\Cϡ��x�n��q��cRqRm_G��'eGg����h���v#��ǣԱ�m�瀎|Z,'�e�m<D(]�KU�������-~!��2+}��I2��,����+~����%�n�Ig�r���9�e���AWsc��"E��+b����f5��;-��]��f�Zt���p����}�J �������Z��m2!`�7n'�d)����K�q�U�N�{��P���^m.m�j޹��Wf�����hP�;��گ��,K��+Өl��1׀�mOˁ�
c<�*�����}�R�0�#��nԦ��'����̧s�F�#T>��,�Rte�3�V�em�9M�b�� �Y �����g�[��^:��R�T�������g͒���.���F-��e�Z3juFa�	ଜa�>�
�ںC4,&�h��f���׋h1�<��u��h��u�V��\���P]�&î��Q5�w!-�}�E����W
d��('0' R�F��/_o�*B{��F�2��QV��Xƿ��I�t��ӫ�p�O�c2�^!�Z�2�&�!}�����������w,*�p�����^\�k՛�To2+@���ܨ���Qh�D�T˳�Sy�m	D�������lK�#�ԛ�r������b$ɼ���2��6�/(e���ޛEz6B�ӟ��a�v3�O�;�6�ft+leFOEM6O����S3�U���4�6�a�?��E-KT΄�׿��r�Γ��҅��
I^��O쭔Q�,�>�סB��X�=2"��\qA��"�CPO�����x.'���^j��V-�@�ƒR�hx�G5�R��!�9A���N��H)^�U���Ux�S@zb��B�� ����,*���+p/�Pt���\.�9�����@[/�'��]���k�:�ęD �nZ����)�[�O�����K5O�ШG���?���°߳�j�����+��Y������ڨ�6�|����:�2�u��_��QN���^_hHhz6n윖��y��6Ssp6G�#P�żn��.Q+-Ӿ(�|&�LĢ��r�� VK���r����O��/�^)1��\���[;G}��YE�w
���$�����z"�*�B�~6��0��[ �r���S�.$*��_��sN���-V f��M;�SZ"k���O[m�Κ9L �����\�Z
[:���N��?���	gj�C��6H:Z�����S��6"�e�2�8�.<П� �N�6��:a⪐*�*e�9{9���R�MSvh8�,) ��IX$�;��ݨ�n7�8n�����~����j�O\_�(I[����0hä)Ҹ��tug��5�C=tԔ~M������q�Ocd2��x�3Àcr�Hg�7I�޺����p3�uԣ51f��ʎ�[�(��Kx��:�E�j��@���T�����s�cŐ����(׼���xP���	Jh�Z�0�h�t1��w��[|�(�A�E�!��tH���A�<7B�=��c�Dhq-@����T��6�Zu��G5[�K�����EB3��t`�z�۝i�e�?1N�f"�l���Y�A�O3{�,���@,�_J�$v�.����f������X��O<[�� ��������<-��P<���Z��A8���d�H2h�(9�Yv�p��*�Aa�e��2A�V�\��6R���@@�=���,�(��2>�{�&�sN�U��|p�_.ʞ�.H�_�OiK[(��H,����Z����4W�b�*�ɍS����C��y�D,��6 W-~)�p0��ق�����;4��7�DuJ�hggr��*q|�@��K�c�u2��u�;o`�h�ʒ\����,2Ru�ok�{:I�0V�����#{���"L���'�泾2��Gc�z�J���O�ѐA�u�b�x�dG@D���֊��S�m�"�#^ƨ��]Al@���M&9x�G�ۂ��ɕu��1}�v�e�������VQ�4�2-}�4��v���K�T��/�r�_L�{G��eH���[�|�@B�@{jh̛қl��2%i��U\��ն~�_�_��*�X�k;��ͅ�ȏ%��VLk�^������1)�8�E������h�,@����Z#V ���T���2"~= �}	Ez��F���;$�3P�D4N��H���#Q��7�DLA��*ȯ�l��ja�u�GL����(���b��te�p��f��#�QP���8��&9ߒ���h���5H@�F)��繇[���]Dq<!��C_���z��>�������ZDa�f��J^���_-m��7�k�Gb�vœ�1�����jyQ�>�M�n����H�n�bX�`�A�vzGW*�Ca��X���Kdp��������V�H$H�D��s�K�v��|�:�R�S�K|�Rzq��K����v
6G��o�����bP���/�X��uטN淅LTP\!>��#U]�uSŤ���~�����rg�g���b	�`Z�~*jr�d�W��4t#��5#�h�8֍㉎o�I�����3u��C`u��g�:��z����V���PA�~{^�NYg��sm�-�M>�^Y"�Ϙ�V7��26������R�ϩ�`b�5H�X�F<�h�%�c��(`x���fc���(W@��Qzg>2M@`�x�x�����n޿]
��q�14��s���,B8��Ҹˁ�G2 �Ve�$o�)�́uߕ+h��W�Vo�����Kۆ��I���)~��?"��o�e��	�J2oɎj[�R\F?�}���g.|x<n��`�v6�ǂ�41�%ImkM�̐O/it�챥����}Hk%pt��<�^�u���X6�4�s���y���F�d�㈨AE&ޱa�s%^Z~����.���Ik>V��7ݷR�� 9�#ŧ��0=c��2k�SYƤ��[��-O�\���b(>��	6H4�X�[�9C��c�鎖~.c�����"`��D�~u�6!F\�g2C(X�YG�-���!�U0gB4�����K¦~��p�@�gL�plȻ�z����D7"�oB�ʈ�U�?���Jﰽ�*��yiM�>M�32��?��6b	iG��rS<b�����}3�c�K;�<A�|+ƹgkr�Zyų�{��Fa�[��s2�fƔÎ�}*O��.�\mU*�j��}:��Сp_�(ywC�OfQ3V�MK���k�o�Q�dܙq;$��v��Ex�F�$�H�p�^^��u*�ƥ�1�߆3o�)<\�HxjUy*�0���V�q���!j��[��ʰ<�.�tg�8@�KsjX���y�=����9���V���<T�-���%6v��
���P��r�e3h�n�s59?7��������
��{q�;����覈��Oѵ�_��Ħ~h$��g$�_Q��!cC��Kv��F	�r�a���a�	��T'��mU��i3���.�wؤ��ѵ;����h:���B'����L����ۂ���6j��?|`Ɗ�F�y��eH�ZX�,)�Z]���Ë]\��H]L��"�V��������8%v��,�"V�Qk�=%f�����!�{Z�"��=�A�	�ml��rK��B���4��/�&(9�1���V\���z��H҄��(:mPM�N�լ�h�M�݄|T�ۼ�9p�s���<���EW������h＄������R�@a%I�I�YIY;$BWYb��-NP�ߢ9��e� xh�*f�]�[$#WnZ��S�x��H�����T^8�B/IsS��2^b���#ZϠ�<U`�AoD"���T@ܗ�[D᠛�!U(�p{\X���|ل�wPX֖O��EE+|4N��a��+�\G9(����!X��n���ކ�$��I�G��������-�թN��f���ȫs׌��N�H#�!kvB����#��ߋ�CsT�����*)g�����&`5^5[̒��8��y�iT�s�����ߤ���"�����ӄ$4n7#�M�b���+@֓$d�I�5�u�K����5����
pf�!�2B?�6�G�R�r��%
���tKif6=�V�V(���z�ͦe٦r:��9&_�O��
7���Z|��`���@/�.�^�6�-�����h��St�I	�"k;&�ɮ'\�6�P��O��]�N4O�#�d5��$]U�Ii�N���X�Nd�Ub�S?�wzP��p�s�Պd�r����/1r���jݴ�j,�k��OE�)�2�T)��N�I&d���A5���B�s�X?�{�%hq� Gp{ ǥ��~��&������Zih=^ij�okKg���c��V/�.��T�葟g�Ӌ/���h[��0iU�����j�f���E��Ȼ��|U]�/��R[�`3!�+8k`���(V���t��֩�R�*>�o�K��n���ծ�Ia�������� ����V�O�䧆!����>؅;aW�{��:w	�eH��X_.���Z��0�t��m��e��;%ZO# ��p��;��l�|���I��!��˻�� b�����mW<	����7O�2Vm�P&�J�`+��S�L�3��r+��G��];�xȁbJ:;VϽ��y�����~P���tY5����k��J� 0?Z�"+2&�w^�7�H��(1�7���GvY�-u��j��X�BXG#|���cʢ!rG��'�ђohN�W��^tg�>�� �S �!b+��!/�T鉖P��G�9:������v�\�řJ��]tll�/�z"+�r׸���M��0�I\S.�\,����f��?m�O���:U�:��/#��ڜ.!��g'������������q���I�>M&���gP �@��ݣ#	�ؕ�_A?e1w�QO�I
�o��&�t��]��]�����]�t�����O�W�^��c�m}+J)u~ x���
�cY2�W&�I�a��������:��+����7c��/5�{�P������� �o]�(�7�9��&O�|[��6��0Ɍ��6��Eg_�f���H�4 ��������f�tK��UjPy�Y��7��a�y���0�����|/��L�w��E�.Бה�4�
��SH��O�'#� �ιS��R
�(O����د��ZL��Ck�č��2b���:A��檸00:A������ݿ�� ��L�]�Z<_~#�H����ᷥ��c��VzE���� �.2I���e�(�+h��)�k���r�E�TW��S�*��X�Ss~��	�sO����Ҍ��N���.*���{\�bx0F�|���:2��q�DQ�>�! ��y���#C�=���x\�'�f���_��������c��P.�SiN�i7[�_F�k��#�#˹�ot��(i���U�	_���\�J�oo.k��A-��Z�%����� ���w��7M�(��{�(h)�T����ת�3ч�"3�&��2�Ģ����OsdGC��|l��S�"^�/q8X�:�|(�u����ujB�O>J�$L��R�p����Y�OO{�y��k��
5�܊�NJ�T(l�r�A�@����Ke7rŦC:W>m�M� �7��L^]���ɖ��H?۶���g&>6�2�S����Q���n�}����8_Y�j�yTƚ}��=�df��*�JveV�R��Ph؍�6J�q��yg�����@g���5�2����br&!g�L S.�5�>�u�ݿ��V�����$�_+�.d���p�����٪�<[<[�,�T�4��. �1��rk?;	�	(�lffJ���_�(�V�vfj�F	J��a��c��y%�L-Ɉx;a1l��Bc���ӻT[�'5���g��,�#t;�����h
���G\)���*���9�4P-k��>�^�Z�)����M���r��0��5�y# ���$����Rw�W$*��L.�AZ�9u��*}��9\\�;d�����Ep��R���a-yz�B WH�٪�Ȉ�x�����(#���w�=F����I`Z`c�کU �x�R9�$o��4[�U�	�&��U���c��\���J���������a7.�2�L'�·iY�8�2���=�'
�li��Ş�Lyw`��N��3���g����j�|pS���;H,�hS��~Zq��}�WOѕ�����?:�wfJ��{�U����ML��s���`5"�*zW�hE����saNe3�-8�5�Bc�X_�m�7sǄ�H��G9�/��f�#�s��>�P���G�vbXr��0��!�^^.���
�^IMc�ܗE:hN�,�}ܼ1$E[';F��J�q�")�Ra����e*s�*��z��?M:ږ�sw���(@]o�M�w��P����4G�|��-a�UhF֏�0_�43�C�X~j{kV :ѷ�jxs/"h��ʈ��Yp5:�ۖ�i����L@3ܟ�h�ň`��jq��h���.�c"�ɃZ��gG�ja�~��k Z�5Kﲭn!�}b��L�����*3�j[����N5�6����;�Y<��Rۅ�	�c=֋GQ��󀚶l�1bq���<f�����I�oZ�cҬL2Ծ�+C����׌�t��x���|��E@ki���:��S�����: ����������]����6���$�9�[�b�y�٤�6����#d�k�Kt.�'>0ހ��������z���=nn�z�`�����+/�@�$Xhm7���{sVc���5�J��s��O�IJc�7�����g�ғ�+w8]Q4����j��*8�Gy�@]�b� ~�� ?r�j[�h��gy]ee��5@k�3��.�u?t�P��	3m0Ԕ'�DA�$�'*���=$<I/�0��c(��9��i�Cig3ȪA�������ew����M7���� 5���c����``y���
�&I&�B�)��v��w���&X0��T*�����*[�+�L�Q%�ha����Vv"~_i��0� ����*8B�e&���R�Lr�􊁆g��U`<].'L�A5_ruR��b�E�Z���p;�n -=t:�W�K%;E�Bj��������>����!J���0�!��dZ�eb��t���wF�~b��)�>t�v����1��H%M>h� �JaIO{S�����#b��w�"m��:Sɛ��E��_�Wx�qĈ��)��@�5tfO�1�_Ü��
P[���:gG���t]&k5�?���(DN��F�pPM~��������E.w�x�!�S ����B">����;�[,ڳB_,N����}Ip4�+Ywˍ�$���S=�
 Q@X(��Ɔ�'u�d��d�c8�K����^�FF^P���57G��X䊒)e�����O3U
Ҟ?�!ͣ�O$�9���O<���N`��,�Q���D$���3>��9��Y�����:�h��c��8�j�VY�0X�F>��[�Z�n D�~TU��Rq�,��W�O��e�A�[��X^c�wo��T��ej��S�W�Ӎ�m/�������e���ɟ;t�<^��5��O���Z���_��茝�E�.dk����N����,�3I�>�{  k���ݾ�)6 ����p+�,�o���+���rw��{���D0d��|����Iml?�a��W��Y�|�ɞ�y%��?>���o'����5	YM����9�0,�_��s��G��*�!�~&��Gq]�����f��&�O1�<�(� n'��Zg���nq���㰆� �����S=��g� �%�j-D�hB3��Y�W��.���Yɾ �Z<
�W�#��j9S�!���)�NKS�4�y�sj����F��p�#�,���ԼM�IS���C�������yB�������^
6�7�n�ƑD1=�M����9ďᷲ�b���៓�m�z�K`D0�h�M���	!]�4��sb���V�q��t�e�>�2�W{�s�>�q��H�V�j�#���K�̻�l�<ิ���ͭwc&�l���ھO�6��8t��R�.�]���^طj��E_�իQѹ|(���F
`#�.Mײ��ISoϟn/.<�Nh�=��^U{��C�k�w��Mh�c��O��������6ת�m��d�gl���+��n�Ɩ�����<����<�������Rp定�. �p]�(^�=��D�Rh<�$��r���f��/M������tF�ǡ��.���%��𬚎��_~�`OFG�Y��^�f)�����`�h�,I�����*����*0����r��(��<���T}+_���~�L[��*u�)#�p�Dj,
0+��X\�m�L~���A�I��~��+�eBHa�[�B��V�]殺���-=�-�)fy��]��9yw�[�e�c����'u?�;H�����@&���
�'yp��	2?6�ֳ�l㵒wI���"�ݰ踞�V%r�$׬��7d[�F`4��7����T(���,2���ކ�ŘN�)�/�pE'}gs=C���L:�.�e���3�s3��f5����A{1��e�i���#�VL%�{e���/KLV%��9�%�3gڲ���O��j�����6�i��>��c�2��C�bDq�9���JMx꬛�q�>�ۙM���6Հ��&E���yF%%����@3rZ�YB2��d�#g빭2	c' ��*7�Ut�h@�ޥN�!:m%~ʮ��9��zȍ�,����p<�R�8ŵT�2d�)��`
[)s�&8�\��8��l�[C)4l~,���Iaʘ8�q�e�7���
W3��T�㌔��ϩ��w�ۍo�#f��j�m̕撲'�W��n�[���$�*�i�<Á��(��_i]j[��y)����OI�^��W�'v�S���l�Ɗ��p4&�m)�X_A�G8մ����*��.��*~;d"+��`B"�N���T���+�ݒ�XoV�^��1|�E*7~�`�Yng��W�n8��o, �bv��[�,��B��0����
ã�j��D���dZU�����s���U�*�U��C��mu�:�- �Ƿ$�}2�[*a=0WM݂o��(>�lCP���.��#�WA5���Gr�\�V���u[�Zb��t� ��9��?ͩ,z� ��,W����-e�cg�줹��n��}/���b���}g�_h�v
c������)�߄l ��}8,a��ްi��I��4	]y��z)�i�o�N��ψ�]oo�~r���-� �>a�W� >��G��7�(�(F�3-1��ݯ���Y��Y�qM����؉� +�Mn�����tJ�� �� �%���Ȏ�u	�Y^����)HBH�5%��B��l���OcyK�)�VR	5���'"���}�W���Xt�q[����p�Q�0Ań����w!�����y�⇠C"���H�����%*jv./V������)� ]���2㴴
��w�B��Ln'��lP�z�ڙ-|ufBF|���G*}Ѳث�4���N�0
=1Ѡ��˚�z��c����'��M�i��k�S��[��P�H�Ѯ�?�I�f*%�.�n��G��Ҙ����WU�
��⁆I=/�[���.��0=Z ٍ�Q~^r4
�2},[Uc�׸���,t��1���v�}� F(���mVZ�5��(�J�e����lL�E�9��D��v
���ֹT �oŌM��(C��~���lQ.I������;�I �~�\
y ����y��~�2�4;���&1�ک`�TNH�c�K�/ӛގm�����=��%	/q������x��:��Q�j�@L�d�Q�)01��i0��͖:[Y�9�bR���}���� Й(
 ���)yhiT+"K 3~���3T�&Pw����:���{V��"仇I>Gz�h���q��{ƭ���#���$���M�z��5Z�1c! ��-?�ܾ�\}c�擄'��k�h�d�ET���V���[�; ��htW1��~��E���k�!�����l�<�j�5D�k�[	ܴydF�*9�ƠK1
�"��K�Jy��d�4��zx�֨V�d#�B��}%�䄖��-{�C�t�]�S8�Y- �\j*�����+�.��-@�7�Щ1�{ș^��iĳh��G�g�q��9���o7�*'��t���l�%�TjxNR��*`�U:=�M���WL�Tnl�Yg}H��
%F㓅yS]y���PH���%�@|;:&�n_�u����ͅ�m I��=m��Cҫ�E^[5��UW��<��b���(��0����/y<�s]��@<i)4���3lgu�߿��?�z�G�������C����澻gb���ػ�0h��Ӕ�)T�x��ҷ�|���P��?�y�'5��7IE.*���<�Bt�>�W*n��9қ�C�]��2�H\���b�%��Uߊ�M�ݼ-6tCaul"�%�)m�ڵ��c����A�t^��AL�4K���]�4}�r�Vv;Z�QN���������Gl��LǢ�4���D�+�/��t41
C�?����j�SP ƉU�\�
~(L\|��3����h)��οR���YF`���|C�yJ�8��tQ�������������F��G'�ڇ���~��L�Ȅ ��%�s�b������nC�St��'�	W�-�m� �MO_;A`�����r�H�o����.��R�L�z/�����D���yXB;آ�z�;�? o
"���d��w�>uX�`n�(��$<OFe����!5X��~RL��6�f��Q2�:F�{��bD�Ž8i9x�w���ٍ�˝�!2ju7Nb�gy(�8z�TDM=j�����ީ2t7�q��jF���p�_�<�;��K�# 1�P�D�]2Z-�&[N� ���Ɔ����� �U(����T~v�q`��$~s��J�}Se�&�ݴ��1N./r�R�Ϋ���1T3�=����7'<��0��R�b�W
X��&�^�w#�L����j�N8�y�&϶������G�Ug̛%W�&�c��#Hܠ�y�=so�d��N�1��Q. кr'���m�u�����·�p�%0�x��J�Iii�����k�9��n��p��j+!.�Hl�]�*��)��
���[���-�/�l_`�r�]|�G���\�'���^�=��ͬ� 2��4_^e����A�H�/���,Ƚw��Az�c�%W:�8�������ͥ���G@1M�`��o�r��UM�c<b���������}N<�a�[�nK;!r鳟l��6�lh\/��0��W�=zf܆~���n��O#+o��� u-7�/��D敱XF��=j�%��m�k^��H���7
)��4���O3_�$�%�0�ZUFM�� ����f��J�~�iK��ad����lT��at�i��H��Z(���fru9\Ш�q�Cs�>@t8m���V+����6$��O��T'��'�K���f6Mx���H��&��׾3d�ȗS�䟢��j\�Ʌ]��Q���r�ubS��"-��f��uv�\QJ��켙�����5�|qֈ�6p�Ǿ=ЋM��E_�2�_��?��NeNJ�r\�l��K�y�&O�%��E �.��v��B	��k�����nK���_m�7:�ȝ�lUٔl({`+3g����	�C��E�}�&^ʮ�'�k���Y�h�i����Ed�uU��������|��9�>����\��d��� ��R�
��ȱ�U�i.	�ݡB.�ū�Sae%�|�s^M��i^��[�pzN-�_�@���c�XÇ��zr�e�K�Bq<m�WLz����v���Ü2�G�����yS^���τd/+�Te����f-/>7�ga��Ԏ׹w?fX{��k�P7.�Bf�,%̣�i9T7�~G"e�>���Ekz��^cT��9Q��qy��k��-���?RG`�c��8Smx�Z�WG����J{���j�?���8t�L]�^.�`B[�rΣ�?��w�eZ��S�H-���?�8^h[�Z�Y�z&�d�h����[���#���%���V�ggaD��.��j�j��~��5���L]e�Y�����@�b�Ƌ�R�?�pq��]�#=�K'�V��KɌ#�)<�7#�J��]��Zd�Y�64�~�Fp�{U��dWPjH�-=�����֯���4��/$���aο����eIζ2P
p1~F^p}NN�c���@����`��"SnZ��=���e��1�^�ӈu�N�K�a���,G��'�%�M��3B��^���"��	�����=�m'<ߤѸ�<�,�NP���:�C>{�PHb1��;ܕ�[��9�]��o@T������zM�9��
k��Њ�0v1X�^�6&>�l]7_�AZ�ߗ���I83��d⭊��(�*)�~��Y��u3���k+S����B0��K
~�,���a�I;iC��BP�9��Wf���
�nΜ�$s���7�%��p 0���0.�;!K9ȡ]n(��_ўh����8�n\l�$K.�ɞ=�;X�'�,^��ڌl"�Ŵ8�)��:����⎴�ɵ
C�ߡ	#�I�u���(�"�9rح\6��t�&n����PDW�C�0��W"�BaU�kB��w�`dn���<l@ֿh�2��L{h3�X��G��Kyg
@76<��Z���DQ���UX�	�J����Gݱ���km�y�`���6�m܁��Iծ�#.�ɩ��c�d��'�Jh^C�.ok�O�f!����r�[�y��YM�*g��-�ΰч�J�G���ϩ�;�~2dx�]F�Bi�$����׵���Ʉ���j�P�	�'|Qa��	v��6S�GrT���|�J6�T�M�\GN�-<B��SR`؃�$ְ���KPS��Y4���㜐J���(��l��p��hsI��⵳���y"j���V?���}]���M�tB��}�I�o�X�ŮZK2
q���#Յ�}b�L!H�ʽz�V��1g{�����OG���_�.�<V�M�Q����Q�y����+@������A�y�{I�N�K�"`q��W	D�qR_Nm؃�P�iǬu��Lv~ޅ���%��z��,�y��>��?��k�7��\ȫ)����$�żb!<L꥛I��}��-�IP�WV�α�d^�F�^a�P&-4���wj�n57��2�=r�ˎo,�ޡ��|E[7/�����X��P;�s�D2Ц�D�� [(��%Ό?+��X�!ڳ=��?�r��ބ����Mt$l�{����+[g������A��7c)�̞}Q�]����x�����8{ޜR�˱֮(���c��^�-	MZ��Aɐ��D*�4����dV���%�2+�����-eFL��O� ���s���Yw5�d����û\�a�����x�� W��'ٲz��n RN p#9d�f�u���H�� G��i�e!<=�e�18�4dРFw&ź���"�� ��e���Hr:�lM�Q���b�#���+�e�|1Q+��D�~�dc�R�f�%T,d��9��}�D8�J��x�G�Ű�axK�N0=�6�/`L%�$���~�'ߖ����B�]�ِ�L'#���;	m�K��eW���"/x�VM>�6�kZ�#��3dp�7M<��X����������ײ���#i�� ���1�a�d�ц�a�B���7�س���ڭ;|l�����an%VK{�3��m?�op�M�{t�)~��5���ra�r��8�)��Ö���d*&%��L����3p�6��C"�A��`�,�%#Tt*x��Z�Z���������� �i[`�%���]�l��x�J�LC�'��l�_e�"��)�OV����=��=r�#B��%["���38�X*�#/�����JL��tg*��LR���U�҃�������h��Y�:�!d)�T/@*�6g�Lﵱ�:$�K��HP)Gul)�R�=-�h��^��j�K�8���q�^��u�۾ۧg��c�@�F:���=)��k�,��@Oi,�5xϘ�d����l�Z� �T�gׅ&�V�������\�[
��Y>��#�Z�%����,���J���]��vM�gД�:�NEx�,-���A3pzL�LS����v�c㮮q�G0���͹�ￏ%�V�$HF:�����!"vYT*b�e�7G�܎=�J���?�.�k�`�F�&�/.��ӡ<WCR3��MHɷ�������� ̃�Y�-�B��A���i��d����aET�"���T4Y�]�85D:���K���M oK`h>`�zB`d��wwN�r{+aVk]�d��V$���0F�%����i'?T�z�w9�F�q ����p������PER��ɫ��.��y�Ϧ�zڝ�x��m�!�Z`� ��OI2�n�P��>Cnk�����(Iy�ăBO�` "�L�!�C�;Ot����T��/źA�(Ri)ۻ��^��#��?ۍ��%�8�Z6u��Ձl�mS#Y��yы΅�������$v�#�44D��;h+��gz1ǳ$�g�'��x[�o@��v���d#�W���(��F8���k���6uğ���M�+F�	0���R̤����'զ�%D�6K�=��fv������:�V�[=�� ��1�� �l0�R�if�A�[\g������8t�b�_�5�.4P���YX��:��!�j~	��^3U�����G}��j!O���nTg�S=��'Gk���g��CLf/����r~���8���N�ׅ�?�S\�W��]��[P͕�����0����wn烠8� ������su�=�Յ�~鰧�HHb���C�t{��d�D�l�+�_�ю�/ԧ���_�_�]P�(�u^#*}Y�D#�uMRW9ݷ�v����Ǫ(�t
���
/ݨM���D��%K�Gg�&�yL�.�/�{�;*z��8u�d�E�C����UK���RsJ���v�|�~����+���Z��m�u�+O�Sd��6輁~h�7t/�78/|M�w/����ˣ{ Z�h�ʋ%n��T���!��Y�^*��!���"�l�B�X[�3���\D��+�᷄5���tY��G�n�[��̣%:y�(ul?gQ�(L�csn�-ZA�-��3�l�;�.�v�4��[|�)VL��͍�%p2ߜ��*�#�tCo��!B.0���_P �;Hq�;�@sa�1߅�?���K�$3!�KC���R's�$��5o&�EA�{��:��{�B5��T%]��*Fp��v� ���������9Xd�E<�����)�<�F�1�1T�BP[��a]�
���	�(����9l��-	,���m���<~����`�����A���� �*��B3V�	<&��4����\��R�O��A$��'_z\��W����;�%�
pMmx=���v$���bc���/�]�S��ɼgZP�|�x){ş��Yx�4-Oj��c66z�A����y���8���F=X��K�^K.^_|Bݙţ���Uk<r���4I8XvSnr�Ǹ�{-���:��/dR1����I�Mb�V�Pf�k��y�V�����Bx�D߽���L��P�Z�Mt���c��vG��f!e����}�{��R�Gf(�K��.��F���?���m* �SFM��E��c�(��$.���U#�j3�`�9Y��I�O�-=^!0K���)��9�2�zZڂF�)��k�����;*��Z�FS9j�%��w����d�5��F1��^�R�N��m�EǴ�������j#L̬��J�Fl��lO��
�
����N��vG^���`�?0�Lq�[���v9���oZ/#���V��_�{����|���5Z�8���0���=!Ym�ɀ�� :V��uO��<ᙃ[�,��%}�*����m���>!}��h�ھ������۠[A����C�����|�"?��!qf���M��fɻA�)�F������tߍX��wzV�vA�y��7�uOR�b_����\�� 8W�J�Y�SZ�W����b@�S������2AD/��У9O^1��ж��j���{�_o ��	��KuG�{`n1|�|�B���Q7eu����y5ᑄ{z��k���7��	�6#Q�4�l���T�1�i�A�'�ena���c�q.�/K���n�&-�dܽ3�µ<��m6����9*�R綀�0��� {Hф���"+��9j�R���U"�3��K4}M�b%��w��w�ٗ[>O����!�=��X�����H*�|�x�rzRfKD���=CtV�*dq%��t���uO찺Q��z�hr�`&����U�3���du��}�u����j��v')W*{cp�u�������`Z�U-?��F"̃zr+z����+D�7��������	�	�Z3=��5=���fa	=�l� �
���pb��.��)�V
�Tp�;0�$
o˨^8�n�bHm���@�$Y��	�l ��ɘ:>�3n3d�#��6�B>��b�N���
��A:������K�N��j�$���	X�m�N�=�de+=tyxE�Qd�����ⷪ���H4���D!L�ag�ܑ��]�v��G���9%��-��k�y�ۧD'��B\w<������D.�Q��6c�ژ������C��Ba;O�)uF.�;�@8�c��c	�f�ଷ�F 2 ��S!����uSK�2`lV�N�_�^�?�d��%�j�./�mx#N�8&ID��ٜ���%u�����9/����?�j�'"Ĥ!�#4ӹ���F�ц��0��b���(O�e��!�5���~��"����/m�r��/�]�O&�/l�F�gŇ~ ��g0�k��QZ���h<����-��f~���~�]��w�ߋ���M�x���<��`���������D�sT���j%�+��v�UՏ� ��ų��5�`$�����4.1�o�����hK�vJ�s���ٿ}��cg��'��u0��围��-?Fѐ3��j��!��3��a�t���떟g��$�i�p�������IBlދۚk^�-XV߅g`~�A ��v7���|�u&;(sW� '׈�� ��2��Bp!��8$;מ�14}�b�:m(�CA4��� ҞX���:�O��Mg��Z�z�B��:�����w�_.7�l�/���94��� M�	t���z ��-]�Bc�[��-0l`Ӳ������$�%�/ǳ�և�w�#$����j��-PAȧhN�!|�`s�]E�����g:�QD�ы�
ɖb�V��A��";�AT<(!�N��#N:�8bWw�gq	��O�f8���&��h�8���xn���ªT{(����;��7�)���c(x,��\�(���}@��\T�Y���m�g��cB⬀�AHa��ٛ�R�~��t�qw�}[���EJ"<E"�_{����ۀ�� Ή����>��b3��^���1�}Ix7��7��[���fS���?��L�şxd��	P��]��QX�wI,ܼ��̣��C�f�Q��:pex �f(ܖrx�����]Rv�>�0�O����H��pM�{gƲ�
<(}��'_T�����a��̑�RyDs
l��vӆ�u��n�>�v,��;è�8��3w����/�}��8Bj�ӵq
�y�J5����[�מt��ss\pY�����B�`�2y���CP��2�����sk���B{�0�UsG;)4\⹩�� �:n��t\{i�4���1Ts�-i�SѴ ����M�;��~꩕ʹ/<�#��f����z�f��dL�J������1�%���C�J�t�H���������P�(E֟��l��-�[j�L0+dhrI�@�;��ph��>Q}8�;��"��t�>b�l��٪9Z�L=�Fn�	W�H���S��%x�GS�3��b? ���^���T q���{�����^��������S� �:�U�]��U�� �_R,�A�9>���298��CV��w�i%�Xa��椿�/�H�= e.���NT�~hC�k��^+��Y\'gg�'p�F #*�8 �Ʈ�aW��V�~�^O�[�ڕ�Sw�ypP5�o�ة����U;�z�+pg^�4
�t8X���X^i������*��HKS��g1m�Ь�����LU�E���Z��R�t����� �v���Sx[8A���O�)q��R\3��M���c�����E�s�;�"�{��j���"*� ��>!��̤�-���A��x;��(���(�@�X�ח�V}}�)+^"�A���/H��L!�3KJ�	�е���ZS�j�<��P�΁���������.�2Ǆji�^(z%ETO���tY�"*Ce���+.a���=?2͏&���0X�J�E�xR�KY������~���0�*�$o��o������Td9
������Z�-'::�=mA
g	k��F�Qmuj!r�ˏk�������0�h5}�+���m�`
�@	\7|J�:rli#ֽ������@��'�_z�����3*Qj屻��"Q*�¡�I��V3�����_or#��M_�=��V:��x/%����o�<|������e��_���R����s�������3p�۱�g�̚�f��7�m������RVl^'�]�p��E��'8f��W%�k�d_�T�$e"�ν�:�Eh�Պ�c`h�dW�"PY���*��l�(<�a@�U�_���!c�'�h�U��� ��heЭ�>rR���{�H��D^C�D{�E�)/�c�2�M���W����`uƖ5،��]UJ;��j̇"C%����)FbTz!2�b��1��ê����Yn�X$8�wF`;5y�kl04���̾�P��g�X�ڈu�];�k9k3��*�����	���`C�{��wz�Ւ�8�=���GO���^|���B��Gm�F@�J�i��~lĲea� �t���/����x8�Rl�@'�DZ}�Λ~mDC�2Z���Y�#���c{�	-�!^F�P���$f��LW)�lu�X�A�k\�\���8�����cR�:Zr����P#�^Ln ��v�S�M��/���sD-��(�2;%K�d5�5��'I1�q�3��lS��M�C��,h� �۶	ұ	ۯP-!�t*�@�M���y7:?�� S���h;Q��^T�x������sB&�;�V�B�h�H	FՕ���%j	 �*�����h�@�
��\�Ǜb�,� 7��s��t;8�=WNj[۴C�U�\�Y��\U�qE<�%�W��T� )���N,$� �,�ZZk��3����*�.��Qex5rh�&������ɺȳwj\J̦�ݟ�~X�Մr�;��0�=��Q���X������7���1@�2fr�h���0p$�?�5}2���ճ܀�ͦ�ڶm�Z�y+��P��vS�2w.�q^S������Ϫ��E�3і�2`��l1V`�B���B9�����u���N�{�~�/z���'0<rL�V5����I�3q��}�y[4�:lk�����P8�	�����$�u5���[��,[�W;h&2��YH���0} ,��@ E�-hޣ����҈84���m	Sǥ�c�=[˯��H��(�2�Ѥ�ւ�[ڈ��(���k#��驪�$��j��Ә�l�P"<V$�O_^�O�)�*��e�`~Vg#RT]k�����
E�CL5e�`a�\�X�OQI	�!�_�:� �v�Co�?�wy�A���=��fb%���d/6p;J�7��b1ñ�a����R"�?u�x!Qvpdv�E�5H"�!�_��;ʕ�F)����L&���7����vꟼ��H1�P��\�R��D� ��I�B�߉�7���*�R�*�'�J\G���;�?�Ӊ���֚�D�����Ʊ�q|��92c�i��>������wL2���xk��j���J��đa����;�D���FZJy��M��Ƣ��ʅ\Ӯ�L#G2pj����{]�إ9��u�wA�6ӗ���4	Ʃ��1�\�(h,���[#^�9Qr��É'��
U�L�iJ��5���2�ib��ʟW��|��BT�Da2�9u���G��KF��)|�t�s��cpu�v���eu�d,��*��ڱSi~Pt}��W1.���Dn�S�0H�OI4�gH�ã䷊�x�2gc���r�g�2�fĪ��N1`2"����
�_�jU��F$�	�)~{����䊤�YS\vp_Hy�����vZ]I�����fR���=#������R�0E�g.� �u�C.c)w��jo+��`AR����Ҟ)���+f���m�t�)қ��|J�
�iJ�^$K-+RĄh���%�ϵ�gD&��������n'�F���c4�{�t,��- L"���D�������R���=s�~�˲�'�6�4|*��EfL"�t3�Qڢ�U��R�t�>�b��|�P֐E@G���8���q�䮰��3�8|h���ڙ/���G�`�A���ESc<!@Րͥ���܎â ��ۿ:r,]�Ty.�0�s!F1��7��І�7�>�n�i�z�+�=%����go�c�d
d#Q�[����
�����oٗ�)�^�>M4#��3�a��I,���oa�l��*�g��+���v��A&�� Le՜�: 2�W��8��&�/��h(N�X�:����}������jo��zV���W���G�/��"ȼH�>Aş��+P�B���HO���X�n;&rX:WG�L:�)󑃱�#k�s����lO�WG#`ܙ���.��SX*)�����Q{<�)\��!y�U/6ܗp��ĝ4
�,Z�<�d�-�/�i�CR�솄�~F4��j�_ݫ�*,��t961kO��{v�kg�����'&�%�0ʆXw�.z���8�G	���l�yY����C�������a��{ �}�?Z/��ī���q��f��
�ĝ�[V��6�j/z,����c�/N�5��S/�E�1�y XԊ3�J�x���"kc|��eq�UЯ��@-+o��O�??Y]�E�j��`A��Yj.!í��=�e����lv!yg}N��,&[Ԡ���;<o�U;R���7e�d;���Nb!ԉ� G�����Tư�?�\�i�U������j�;��a���Dj3{꣇�K&����G�M��8s��ꁤZ��O�����bO��V�m\6��@��_r�lH"����3�1OH4�cʕ�++�`�
��^���d�o7
��߳���V����#FF�໵��apﶈN@�����RO�"CaȜ˾9xυ�<��,�ˆgUN�Hl�.�<^�@�Ԙ���-]ۡC�W�l�Sa��<H?I5��@�w:�o��)1���Rkl�
��5����c��F�jTa��T�+�Z`T��0��]&�,�L��1f�M��\��bP4H�6�c{�� ����oWb0�"�r[:���x�d"5��YNx+LǼ|�߄+�`3�Yd��ީ�cyU	��N�1��t�mg�]�{�ȪR9�A�!�Cw�][����7Eq��J�>�-=#��X�/��M�J��s�Nf�6�M�i����bIP�^�~�m���Z�Q�N�.��;�͇�5����3�R١��zY�����j�kp�~�Qo�<ɑLVZz��|���Bg�/u{�3��Zh!'Y�WX�t��z��I�J0�u�N�v��oL������sz������I&v�(-A�m�Jo�6���=���Ԯ�]���|Ǟ�ް�d���������������ܣ��*8�Y���ԳK!�'ǮX�5�w�<H�D��l�r����<*�������*��ɿ���3s	D�$tJ�%JM	5Ð$ʇ�N~R��Z�R��S黮���
~��o.��oo��xK��"Y\8vax14�p��>?�^�{��iq�~�a<���~ĝ	k�(����{��4$�vf�g���ć�"?IT���(�C]��6�Ʊ�C��}�_�$y8�PE�DP��ս�b��{�1#k$�r����h|�R=���KN?�s�f����CZ�H)��Vl&�?I���ś${��1�I�3����_����[d��+P�F���s�_*�:�2"������7��/Tl�$���d��d S)y9�dX+	������G���AU�b�Ͼ�R����՟��準O]B�_���6"��+"�AJ��"�0QIjO�S+d����^ͯ-��L�w>aȸ�N�dܢ��j[��A�ܜ�B�h|)�3����W)��r��u��rz�����)����;��|:�n����~��C�#��RD����	���T�b�H��/�G�j��ĵ^d���o�m���\A��K�X��>j�������ɳV��B���N�/�M��94,k�]��Q� �5�5VN���S����O�됭k�2 E$"�?�n��Ed�9�1��9\J��s}� �p��B+@��K��w�&��B�T����.'�Za�L�wìK[7Mw�=p��+�#(sf��?
�����.�x��/�5����Ժ�XHՏ�~�q��|��w*Mk��ЏN.���qw� n�>�>�Y7Z*��߽��x(`��Iᴲ7�;D��kX�D�;�~���2��ZY���Ϧ�e9�h"�
$kG�*�Y�^�˯���B�(ʴ�0z� ��Ʃ�Z�\
����n9�]T2
�"wJ�^�N���3�>j2 �1�X�7tϵ����Ď����_�Z`[�����B�.#g%�4^��9n�����ޭExM�����z��&�NK������X �P��Y��r�"b\��]a��/c�ñ�|��e�B�f��%!�ѭ׾Զ��fPc��*)Ζ����蹬d��Y�Ci�X�Ur`ٗ�?o�mt�9?L��^�q������k/ۋuϋ��l7�i�4�h�P��/U�5�6fIt��� MȺJ(�bA���{�ab˼,��NL�U�wlu�b�Q	ؚ�~m6����!�:a� ێgZi.�o��I)#ԣ���	�O7M%m��z:B���~ �M�,�]
�����/�G�n<��Dk���[�.}+Sׇw�?'���mmn�k�Le��_<��S�\O1�㛦_KD��&�m+o�Wޘ|�!�(�h(�bƨn�Ҕ�RK�p!@��
K�<Nb.�_8�W'���t�'�Pi�?-Cu[v��P@�F��h���&,;Yl��e��tW1���uE�F3ĥp��[`�V�	�he�Dc%�_����!��Q�M��ȘW�!��,Ȟ!�w`�EF�~�
��w06۵���Y]�-����������%��:!���Q�|-jN*�)��<�FrsE{�CMJ�ɱ��E[�D�P.�؁�~�����6�y��d��6�=%�ű"~���Y�֔朜��:ek�W^���R=Tσ�L���h�W��8
�"P��J>����T.r��$`�㳟�myJQ a��ݍ���<�~̃�xf�P�$�BRwY8�:z�������3af''.&�a������ֻ݅jh@��v7(�^��;v�DSZF��a��
�|6�*؟x��7J�4�$lb���nk8�'�X����Ю�)%�q3�1S#j@L���c�P?m���S>���9��ҟ�U�O��Y�Z�RRf�#̆�v��k�WU�ϑ$<n���ORu���k̙��NDr���-X�\�CW�����'9ѼqSkI`���p��8�T?}��? r0�%�����1��'�
=�(�gO�t*
l�}���׳�4���0���*�X���'�2�c���d���0.�~m\�{�VE�҃�ժp�4X_�v��{Fb���mw�>�:��k�d���������y%�iA�Y
��6�3hʰ�"�q�Y�8􈄿%|���:�<�_��@���(��z�W��j7��'�oC�k�U:a2b4���]\O�'---u��
#A���^��?�{�IVb��N�R�y[���A�CLh%�Z�f�E����*c\���-�f��Q��ۭ�̣���3=c��Fg��O�ץM/F v�@}�3��2�{k�dv��lPծ��d�/s�d=��K�-Uc�ZB}O �)hCX��2U[��8G@ �TT�n&"��,AOl��q�1&��O�V���g'k`���r���R%�ɮ�b�^�*��̫أ��SYsZ�<֑���w�Ĵ?�MY�V-u2G���o
u�h'q�_ZT@K�����E�j瞑�WQ������'���A�ش�!���c6��Xi)Z��cx3_7k�p8��$�c-�(0y�?<��^U������k'�6��wj�,X ��OTT���B�;�ü�1ص#��)+�!'6	/^��Kl̖��@u�^eG��ogm���(�z��N6���"Η���R?���"�T۾��@���&��q|�^�>'�u�ޮ�,�e�D�i�a�#CI�U�3��%�+k��z"������(%��FR�##���L�(�){gj���lTZ�&�(A�� ���4�k�;��X`u3P�$׃G:I5��vӦe���I�3[˸S &�*Ak2�f J��,�{%�~�n�r�D\�d�}�o�CG�Ѹ+����F������gkt[Iޒ|�����bp)�F�wL%E7�[�NC��*ý ��Um�����xB!_v�qmu��.��*�!�Ii��O+#� ńrD�,z��	�l� l���3kn�+���Pk`ł'�2�P=�^IXb-���}�4�4BOv�&�L���+ӹ#�~��C�M��g5$s����O୧�в���+��]@���ZG 5�T,�?��2�RDw Oa���1�Z�����=X*�1S�jY�xyx)�<��=y��%P'K�a��Ej�bظ�!AQ�<��z�L1m��5��]�$Vh�kYe��\S��b�m���o2��8B�@b%+�=g�r�.�4�^B_���[ ������v�@�9�}yp~Scۤ�*�f��ČA�� �C���^���8�(}7š�m$���������C��s�]�
 ��w3�^�I����8���V�h�m5F�VϚh� �K,q�,Ę���q�gRi�i+R��Е�<�������I��<��Ӵ��K��q��	l�2����p��y�$-�o���v����S�B�7���S���ö����V�!gvY,�?�}��l���w�T=o�q�"=
����¬��zW�O����·dM��8O~7ǵ�?#�s8Y���s!zc_�gx�:8A�������ڊ����wts(l�M���v��.~�U��S�u�#�;�-��V�5�i�w������q^w��ِ�qP��Hn-��i7�ޔ���qʉ6��=4]������X6�$�8
��K����t즧���z�>$���*��������tx��b��y�<�!f�#�QJ�F��8 {�yu�^>��?S��	�e���r=&�l
����J���.��P= ���"pY��ڜ8�ʩ�i��ڤ��eP�xc�;�*�p�&q�?�d�# f��ܙ�������ue<C� i�?����˸V0È��aY�N��
�#!�*a�(/��:~���vp8��1>{X1w#��z�k�:�R��UD�O`��h@�=����
v���bv���c������g���sj6�Y�.q�mתkX?+=#�\*��8/���������F*�~�$����&J������J���;��-=(я�U�d�szu��xr��ۜcd�O�֡��<<�r�F����,V����u����VM��)��"����ZZ؂��<}��n�c+��H��9<�LF�����kbW;�+���e�=y�*�ɔO��%�H�H��<3�#�����R�O��*Q��c�>]������k�JA}*��#Q��{s�]D�]�iN<���f�3���h����S�E���r׻�y��ʈ�1#w����cW_o5yN�Q����b��\���/kag"?�<���KqH�A'=�ypxU�Vo�c����l!F\O*&�����#uc��O�	bh���Tfn���5��H�,�,�-o��$J�Ce�p}�����F��e~�}���צn��! �J���6�<Ѣ�Nw ���z�u7��;'�kq��೜ugP�㬦&�η��l�ҝ��4xh�I�Ҟ�Y�%�!�M#�0��E�%��X6ci�o�qx_�
�X�ԕ���}e�$���|��-Wo���Jvs,}~�cV�����r�r����ȿ�G�W,9��Ӹ!���?LtL1�.��h���̵R(o6�E`�"4��-� dc������"��2R�. \��&���&A垌?S�e"���Vf�U���7��5G�@�`*��}���-�ُ�:(P���&� q�c��b<YHF�P�ǲZ� G-+�2DܑѩA�o����A����;>���}xe�1�{.���tab�u��
��|�����߻�M�R��p��z�"����c��ڍ�'3��T�՞P��Gv̔�]����X^�
�f �r9��s[u�����|�Z@�~\�n���N��2���{��8��YZ��gHԗ����H�� ᰆ6-������,73��J�ҫ+�ћtCD��B[���U!��ug�z�/��Ma�]�������� d����n�K����玕��D�E��'M���' UUǕ���:v�^qЪ�4�<JŠޝ�ˎ5M6f�[�����{�w��7,�&T�r�۾�SrKj�� &X$.VE@��u�IRm��j������s�쾢C\�pq	�wa&����s� ��V�"0�P��E�W���*S\�(��JG�5Z,i�m�w\���1{�F�������ȭ�'g�|�tQ��0��['eeQ&���u��Z�g��CӍ'2�T ������-&R�
�iu��p\v1�Փ0������^�5C�:o�?5�����a*{�eŬDn�N��He~��L-.%@ã��t:��C�BI�"���&)��������%������"��F`c�J�G����weO�|"q5L`��z�%�#��9�d�71���H��W�t�c�h��.-���Y����Tb{��3��=��������j�o�\ܶ�0R����|!�[sK���}$#0��f��L2 �u�i%֌�j����ůx���#4���=��8GJ�I��{9��Г�q8-����{��~u���0��/���0��!ߠLZ	���R�������c w�K��?�^kBn�D�kǅ�C33.s)�����Nf�	�����iG�L���O�ߪWW�țp�ERD��ۛ	�h���j�66[.I��~ހ����p���eD��>��w��M��A�������i]�b�����\���`�V�@@!P�����rR�������ހm�+���_�gH�d������΃�-�X�T�U#V/a�]]8��$�%���f�w��pFK^ *�R�"g�_��\Qd�����^a9�k���

�T�9����pcȗ�#!�V@�0�O�M�>��I�ͩ4�`�˻�,j\A_G�콳�� I��>�8ߕ	��Ľ�.~t6s	��{R�,I��:�~���O��pj�Ώ��1��Z{��ǥb\��Y�-��dM���br������ ^3��	���f�S�D2ی<� �p�g��0/�j���� �	�4	���d@/�p%M��V�tFS�O	�3#�-.�e��[4)>��o��%�FZ��:�?#��}K����T�d�U%�'�=Q�) �o��T���:YuZc�!Nv~`5�·<ʴ�Ќ?�cO=�C���D�,"Q�a����?��[���ک�};tѽ������tZ9�f)^VWY�FfxY��8jf�� ����#�m���A��v/�e��;C�#-| ��=���3p2�&�z�a�W����;=���F<��tƷ׻��/{�����	D1O��%�"��Ѝc=�*��wW�ߕj#� ��h.JB�R/1=$�</�i�����k�)t�M������,�y�K�~?#�{���O;��w�E���\�:�O��}���*��"����@J�C5,���<�@8�@.��"��l�O���$�P99�����.���d0HN����jkXq�޺�=c�����/�+턂�a8!adE��X*�%L3����i���^��hh;�f%ơ���T�i)�^}U �8v�"4@\J��D5�?��'wl.��u�q4lFd�ςֳe�ޓ�k6�4��X��`��������
xa�XР|�P7���X���g���(\��uq���)^5f�јcB�Й�W˓�g9� ]�fA�,��ڱpL���ZAz;����$�T��*S#3U+���I0G�O������>��ra.�Q��v��	G���`�ܕ�,ȧ��'��E�]��7�&������'�7�l{�+`�0�Ӣ����)hvf��[(`
�)���O��x��a�� �Sx�ku�%��l��������Z&�Ʊ/�n�Fa���!��d��WKX^Zݢ��R~1�F&㱹l�2�F3�wɁ�y��G�pq hX�����"G����{j_E��c@Ó�rkv+< �Og�<o^�]���Ϙ���=�|�t��k� �\�<w���nß�D$aG��}蟛
{ރ׳�%lޅ��$pa���2���\�Q��cG1�[�~�	������'�֣��w��w�e�L܈�a�Sx��~�o�s&@�Z^o5u�?�����f�P��г�u`.���J��˧���������'3O�j��몇�lf��kl\���;�sJ�i�>�m�íV��k�Pa����d5�%��D�I�k��0���=��.W��h�!0���e!l���Eh���8���G�`�4�ZWG�sr����a�%um��ۄ�y(%ԡ��� o�Z�1[1�$����H�K��M�;[�5�rR˨�|���m� �\�+`N�*��������{��n�<�����Bz;����Ef��9(�R��H�j�h���O����B:�d�_�e�C4V�k������b��z�����Ӑ��;z������ϖ�9�ý<�:��ғ��|
�����k:���
��i⥂^�Êz�n�X�&�2^�fU%l3"޲l��cei�//�%] /�����l�_WW���z��:l��h���Z�U�ʷ�َ�V��t��^S�i3f;�+E���;9���'�QU�5 U�!ĴS�/),pA�0%�L$_#�K�-�ʧ@���`�l�v�,��0?��Cd���o�L������a9?����b�	����#��KL߻X<����x�tBx�8V�H��D��b`JӠ%��I^:j�������*��qe��ST�RtI�@�:�:2��LO�Ѽ+!j�4"H�7�h��z/�!J�e\���e�r�F�X+1}_�->FGX�"�ՙ�{Y���G���rL_��Z͟�ե���N���`��zd�.;VUy�,XW�+�*��4�D~p��E �/�bl2�2��Ikc�27ORpp?�p�S&d y��m�vP��6����xX���P:�|8-�ч�{%�M�:�hߩA�ҧ���̉���D|�º��]�������l�*DCrD6y|{�����ߕ��W�"th�͢b��f{3�ࢤD�R^�����x{�ұAG#����޹��|����[��k'�L��5d��}�8N��t1s��uP1L�+� ���Z]�`�,��F'f��ȶ�a������-��O^�m��1-E�d$Q.��>�|��$w9e�&5 lR$8��b]m��C|�C���<�yߏ)��Ҹ� ��zM���2lGHӮHs��8h��������SP�ٔH���4���_���^7� &cO���$S�Gͺ����y��(3(��<&�m��HZ56Y��Ey8�˕��&Y�RE|�
��pc���CU�v�A�,�4�4���a(�1_Վi@U�[|��3[R7��0�O1�d��O[9"h{U;*��ճ��}�*(��j.��)b�FyP��e�����@��3[�ԣ��!�Z�JRT/�pj�a^�ۣ@;��#��M#U�|���)er���=���Ĝ�ʃ�����Q�d!�ظH��SغSW.�+��/��o�@沚ƪ���Iv��� ��Z����Ha.Y��3_؄���lt�*Rw2;]��S}yC�	¤���8KoX$�i��~Ӿ�u�wHydk�k����Q:���]D�4�S�Gz���񥗁gE���_>�I�7���z�%�ڙ��1���
�O�y�� �(R��N�ѐc�S��F5�<�ᢕC�)�`���LX�2���U���H<�A��wՊ� v)�ɥC������u��}RxTZF���g���܃~�k]���|��m䦚�%.Ǩ��TG���(�3�����턴h0��I/���	�v@�s�0O)a����ל��Ө憋�R������g��	l���=�e����5��T�Ң��T���}�@8���}�Lo2Wp�N(��GLl]���p���%rM�Ո^Axi2]=��.�Wl)z�O>W'�I:���"t\_�!&s�5�S��u�O]I�	!�B�H�T`�i�� bSt�p��	�n������m���c�����i������1���!V\�V`U�X9�@NF$e���^[*b�㐲D����Ұh��+'��V���m�Vd��
J,������s@c�n^�����C���ݒE~�䗽=xW�%&��޸R�<DkRQ�L�_P�I��8�bO栮�G����LF�7��n�-��|O�~'4p��Wj�&| �m�4�6)?c�6���Q���=9��W�o����<��'t�4�"]��h�V���RxMe���x��Wi��l�t�`݉�n����˒Z1�AX��(����5�tx^��읱O6$L���>5s�]����	/9X<e+�p��@�D��~:ץ�܅Y˂��i�JbJ)�� ���JZ�a���@'���߈-*���.��Zʶ�&]{e��Q���/�u8�����pt�4��E]$����~�VjY}�c��&&+7�D�[�+���Iv�[����0Pm�,����ػ$1�����*=��$�^	>ǵ�̷?�hlns3B�S3X��֋1����Ë&����έr7������uJRn����&�l����v+�I�H�r�S�þ���r���]8��u2��/� �]�M�j��#JW���cE9.�ӻ�#@k�2CW�U��U�`��a�>Zg��(���zVӼ`�yY�V�=��­1�y�lM'<�@�c�����|IBw�Tk�����X�zqgn��E�-q�_<Е��s�K.}C�Ӭ�j�D�,��Μ̲bK@�q&��ʴ��] �6������m�v�J�K�N�9M�?�>�q�m�N��i��$ǋ+��"�A|�J��}!�&��.Y�
h�v�����(��b�����ڡ,�?(���I�Rv+�b�pN�V�m�x�	˩2�@�$<�(u�^%�#rk���m�	���?��ϓ���τ�A���z���4j�s�� �VĄ5+�/��.�����o�>��9�M���K�ܝΰ�E�}.bZ�# ���^��ID%ѳ�Q|����|uQqKG���Dk@VĐ�A�ԟǘ("��n`�m��&�Ѓ�,�}�kGTX@�p�iI�*i�t���%v���1�¨��u׎��Ȝ�X��&*Y��$���B��^�I_%'ى�F��"�Sq�UG��Y@��qT쑻������	'��p��EY�j����}SS����,Z垢V�����$�Cp!tX�Lx�� �t���!!��hU��+1bD�9z��ܻ��V~Jwml9�dj�dȏ���&rZcY�i�+�$��32��t��tU����v~�]"������WԈhM% ������xu�����R$p���3�����Qj��_��2?x�R��H�8�]�5
n �V"]>���;-%$��!8%����k�㷸�ُGq+,�_�/�o��H+BM:x*"�R���R`��+!K�2�+諭C���=�vz�Q�mԀ�r.��籟��i�2� P[���dqME\ȇ=���Y��al���E4�8Jz]�i�����s�U�?�˔e�3- �9NIW m(7���Cn�,G���+? H�L��7�k�Tï���������+	��t��ʬ������Z��[b�5l���
�Td�_��k��.2�} �CjLc�C��lXܿ-�J��F]�r,Ч��2e�v8_���d�Z�#��hò)N7e��.Q_1ED�O� �����G����)�Oy/�6T��[2�d��=�i��	�fAJ`�>�W�1��6�0� �.~f�(�����wA��ڟ�e"A�ym���v�Ԯ��/g�;�/_�Vj�-�m~26�v"�3!!H����\B2���F�7������B0�f`,!1�m�s��B�Eۍb�t��7Ȍ�90`���0�q��SD<b��!{\�
��2:��%�����ƴ���-��d�z$gǩ���[T�C�ɴ%-K6������1��͂$�q?t��qRuw�U�R�e����l��O���+f ����.~�IE<������NLU5pN�q��Ƕ����3�E��<��BEb�`�/��G�dC�6�HO��G�z���_�2��^��߼��
d��Ӱ�@LA����?�� 00zH�#� ����BA[��e��Ɠ�J��Bڔ8��vCw[Rh ��J�|=E}��b��f7g���R�F�&#jG�U~����*���h�^�|�Jҋ��g�O�=*p�������LbƲ��v� ��8j0Df�C��v���;�O.�FE8Aq��:rS������)��ݝ㉝�G��CI�[�t%�y�5 <k-��&�.x���=w�A0�݌��h ~I�����s~2�YnԖ�J�C��dN/�+���Е�Lv�dQ����ۧ��r�:�x!s��!,��چ�d������"�Ԙk�{�bhK�g���lp:����gB�>�g(�Ϩ��!+���}���k�sJS0�>O����.I�{��S��	��|c밁�
mWQ
ZD�S7"���f���J����([il��i��xJ��e��62V�4R|�UǶע�d��τ��9�@$��>�!�QY|�D�&��(*U�ev��xg[@2�n��C�#S�p4h�>�ܚ�v_�уJB���٬�8�fwQ.ԗ`��pǘ{&�M���>~�t��Q�R�;�&hC�Mp%�t�x`�h���\���'��Nn��LD�
h�`fl_���#+�7�):������]�a�"��q�c�F/��|�Q�_���ϸ�!aG��#�dUگ�v*4�o���L��	�[�q�?V���|��K=E��[ ,���Z���i��!x�&���A����I%��V��+�x,�����n�r� 릭~g�8*܌���^��&��$�3�NlPG�D�ct��b��^�Z��*ʊ�۲d�� �hR�~�������՞l"תX�Ӗ��-pܟ����m��E�:��9� ���/s��K2z*�)�ׁп&��:�b���zČK�BO��r���t6`2d�7�hH���.���H�Q �xc�ն�ф�kb��q]�$���[ Գ#k
2QԺOC�DK�U���f@��S0��K�mX9��Y��*�۪	[cu�����������e[�z	l�8�����*n��=W�� �h��/�s$xa�`��Y�U����z��=�#��-�#z�כT�8�|�K��X���M9�RHD#e{Zy���e��E#>`.FLa?f��L�	AW;0l�f����Đ둏 _��āi�u�s�*cY�֏�L_�� �X��~]t�%I���}���i�x�'c�Ƶ�g�P��H��P8̦� �&���(�"YO���yڛ�������Ƙfƴ(��1���:C?���K�j��
�q��( _�B�K�~���O)y���S��A4Z�ӛ�T"�P�;ӥ�̕��\L�tdETE*h-S�a0�ϳ.�i-���C6��ߙ��~ϼ��Z
�Z;oҶ�U#j��	��#m�2�@�2�`9h�r1r	������Q_�0��i��؛��AeQ�j�ZC�.�d�`Z�5Z��Y����� ��H���-b�kw�50�O-��s�k&Q���(}��;���E�9D�:k�Oi��d�N���c��~�@�Q^��s�6���ߊ�������W�A*5/"D�d�c��]{���>�.q����(��q��?R�(���N�eB���&��
`Yi���6�[�׷��G�����r�A� r�WT�`�ze�>i��
:#ཉ"�P�O�3|+}��^v��lf�xp��7b.\�A2Pp�����	4����WXD1��p�j�LOP�Q���*�"��x�u��T�c:R}����c|D����4bk I�����J��������/�'�v���,|��ds8>-�)\�q�*����Y%�q%ߊ�8�?0��vC�KK&��Z�
^ �4�R!թ��d_J;�]_ӭ���[��cÞ�cR#^��i������;��<����r��0x�pUx��0�m N�w��/1�ۇ��}���a3��������0�W�Ǥ(j�h�-vL�@��߫_Q��D�(tӺ�Z٩A����y�Q)������!��C"+�xwtG�7OV�c��f���}(dU^[�&Z���t��`�t ��	����f-��$޽����)��Zs��ފ��G
b�DN3f6C���Z�3?���W�멨5�|uLb�R߁F�g�W��q��z,n�W���{��~��Hk2y��\`u��!Mr�M6iK����� $#ƈK�m~���Wz'r���'��i��GqU.�D5���4	��>^=Nl�cȚE�O+ۇ��hֻ�N_��<��H&��]HGk�OeǇ�f��:}��&��?�[1]?���=�]�����y�f	t�����8�1�V�����`[�aC������"��M�<�vX�Gb����������o/jL��Or=F����l�S����c�[H+�\�)�bB�'	��T�k���Ӣ��2.&�eH嵚��	�6y�d�$ԅ��� ��j!������v���S�tj�#�Ab���t�}��p	��kʕ�e7�^��T�#����H�!�ї�AZ�$�i���QE�� ��Q�x� 8*�U�l��e6`�}NϐC�rS��)+�~y�q$����b���hYV�]��_2��H��Y��Ò,�K)���b(ݰ����?4�iX��!���A 8}�3_D����ڸ��H� YH�7?���S�.���l�5�������ܨq:�В�3Sp��TvLf���dO�Y@^�卬�B~�0�ϭ2y�j�{�7�e�3���/?}��ETEO�!3�����!qX+��^�(�r(�ӭ G��4 ���W,2� K˫���n�b=8�ip��Ժ��3x����~[��3�� ����*Ή*ba+|Kx���eEc*q Pu�Pe䥫Y
	�a�s0�	�����PRD����Ϳ楙�������I��j��K����5�y��k�ęwx�)�:�OL���P~���͊�	b��VY8�J��Uy`����P?/^6�w��"a��OdB8w����2�7�d�S��w/��eV���Qӆ��� @g�S�Z9�=Y�~?��K�F{cI��տ��Ϩ7���!�6��&?�����Ê�m:�$���I�[�o�(
d²�����7ˮ��a���<��9c^!�/�<C}�g�֙�2���4��= ���z����P�;m���K���mv���<�`�M�#:T#p��K�z�u�#=M���Xb�錕M����j�V��F���}�=�W�gs��u;�^����u��1��G�~�1HxFCU��9�51����W0���3Z?&�:N�*�/R����*��c��D��l��W��i(+U� !�A�YY�dz�r^�/�.��	���}�S�
���t���"��l����~���%���t����~t�AR�Tl�R���͒�[�0��H]m���Ы�Z�q�.�0�� ��=M���q��Q8G�NG3%�Q�u�X;ח"`R%�����?Tu��!��;��^T4��
0�$��B^B�8QxL���%�WY�pÜ�L�H/�a94�0��L�L��t��0���F'4wh���z\�v!J���KM.^(��O,jG�E�ijsOG7��O�c��Ӕб�*��rO3��j% �3�i���*>ߏB���`���>�p@�, xr��.'�$��|��/��!�l��L���l,���mh��"��r�߽:�~0�]$�up�Z�*���6��9^|����sԊSi4�!~fj��Y߶r"9,P�( ��(U/&���P�b%ΫJ*���4Q.G�ԠE{n�DZ;���'v����Q>�g���E�	}}dA_���&��&a�UN�C��]	rGXG����B�z�½x"��`d<�Ƭ�w����>�� v%�~҉:�g���b��j��9J�d��W��\����3i�2���\��;;�N�u$���FM'�Ծ��gˉ)��q�����slK�ٰ;���Ӣ�ج![�6�x�(m������f�t�m�ȯ�]�b���;��6���k�p~�[��\D�V��ݚS�n�^��]P�{/~�4��~�FVw!8���i4�y(�xȶJnb=X�{����J}��0�Wr����8B���R��K�/���i��m���
ħQ�I$��+yc�ŵ(JЯ�_j��;�)��"�i���u8E�8x�71��n��.�����W~���#�<f;:ϳ~�a�h�M�d�4���+�7<(�81Z��B�l�]�]T�z�O��@@7�$D��0�����v�=��T4�PT
��c�=��6�m�f��ĳŔ�edGAo��[�#a�i0{Q�db�
���d
#�|�6)6�~��]����0X�
��IE�L钉����q3�W��}���=5���O����pc-	s�C�~8��?ez���l�Vu��A��6�� ���*g")6/W��u�sN�5�-}蟜g^o	��?�!\
ҿ��;Q,?��8��TX�����]���Y���'����I�A� T7�	#eDGj���Uy~�� �p�u}	���) ~a��L���#h�����e�8�9I���HK��
sA��R7�c� Zq4���PXvj�"�����O���:!Y�K��mjEh72��/O������(������|�h�/���,���-��WgkU;�Oqvjcȉ���vGp�a:bW�q��w�a�`o�NO�L�1��E�V�?��Hb�>JB+/p	�jjV�冹��EU�jR���Tn��F�p�n�A�nGYC��ZN���hԵ�{�k��8X.�@�4���)���$+����W5M�y0HI�T^o�.=%�;M]_W�5�*a-���Z}H[�ݰAeĝũ�I����`���$]���o|�,F��H=mrdWO�yC6*a�rM�����	���ć� 1e߲�/A�����2I�e�N��ω:��bY?�c�s#������w
0�̡�~u�Rjׅڤ��k���Yㇳ D�̸��-D-��Bͥ:Ձ�������i�@�
SL��Jl��=,M'v_��gMQ��P[ވm�}}����Ҹ$�G�E�]K�"�b��у��M��r@F�X�/�ϊ(���ڻ
ɚ����_�H�}���0-��Al඲�A�#:���]A1�����ib9\L�_�*�<П��7�N�H�Ş���@�r�a] ulhn����ۓ��0e�1�|@O�����W��EL��&ŕ7	xq�Eoq�}�W�M�OX�1v-�ݪ���'��8�����U�\}���Lʙ�$݋��㝕�?�	�\�dW?�qZt�@D��yT��Y�G�~`��<3~��4��X+#���B��J��!�n�f���%Q+N�Bou�V� �	�3���B1����n�ZT중�P��sxb�bFeߔ�+�A��3E�!���
��������qW��m��0'b������ɳ���,�DEm6�O8��x����ĨT�L� �Ϛ��ғ�cL�y�e�=]�!`
�\��M	�?���2+"-�H���ا\���;E
}S�W���׾Fo�m���� ��)�w ��.~j� 1��$��cj��"7��ބS�NA�k���7�1:���-�'���)�l�rd��ڛ6�
�+A6�Zr��樅PrS��N_]�7�r����B�Q���H�����Q�v�D��8��B�;�B�ɪ0{o��z"ە������҆���d��T��&�1)�P&��'��ū	G�������]�!n��`mx�б�4%�ߙt
�,	=��"Ḅ9_]0;��so����iٳ�����1W�g̜���%��Vc:��?~}�f	>OW�Z�;��	L����_�,�:��(�x�*:��d��[H��n>.Q��/t�KI3�Ow��:r>q	X����SE ��ޤg�0�̨�zsh� oww'[�:����'�5}�`J}/��z�;�3]O�����,�AMM׵�Kap-V�t;�t�8,s
{�� 1J'=��-�(q���i$�#v� �O0!tm)ٙC��1�#�����"�t�7D�s1ܣV�,#�Xb�����^�E7�����@�f=���h�[�p��rc��������XP��h����èz�v�O�6��9)s:�� 2�G�b~m���E#7����|hV��jqgz�>u���
���_ì4�J��_M#$���ܜV��#����Kü�h��g	4�����:��mH��"d�����LQ3,��BA�+I�ZwN�cb�p���pC��z��w��l��S��@��˿�������?�p��4n.��y��o"ښ���-:x��wVx�&g\��=8R(4I�:���'�
�C�`oi����#,(�=����EJ|pG�~��I��z^��Ǳ{ռP�`k�����]�`
�[�N�0��M�t^|��M.���#���
5At���ٹ�ơ0ru�hg�^�>�3Ь�X2���#�ǀ��_�LAB_Ґ���n!�ѹ�]�������	���Jj%UF�(��(��0�s�ަɅh =y�@��Z�ն�i��9j�c�L+0f�d�;��0>�P��9�y��-���g ��QI��a�B�֎��#�+��
�z־U�Iۙ��g�"<�b����s`"YA� ^m�MV1�ߎ�^/�0P�B�ۭ)�˩��|����c30g$�3n'�݈�����`3����1�з���&�.&v�uc�y�go����	ڗ�;��/%��/��?��(��F�mL�'�3dE�v��5^��z�xC��Xä]-V"sGg�4���G�#=���l&=
��j`�2�}%[.��"h�4ך�G�g�6�w{�p\��03��P��f�����"�Va�S)���E��Cv�}R�c�r����\��d����-ؿ�HT��:���^.����kaR��r��}EH�f���*V��B�� BzZz�yš[_�;n��u-�N�~*��b��l%Gy�ݨ����C �_M%RE�[ӏf%����k���9\��$B�rS..Xq�Z`m
�86x������9h	�ݾ�>�a�eb!���M"�U*�A8�:uP*��E�����q�����z �.�z�m��xtH��������=�)ef]{>�wՏ�.�q[$Q���k4,K"e��}A�Đ�kz2?�n
�{~Q�|1!tɣ0�c� �<h���W�W���2�����}�.����"����݄��Qn-v�X�����!��+#��|���p��8���ؖ�x���g���"���d�V!i�\��A��N�ϝ{�w�S���)�C ������1O���}��"W�n�R1	�Ъ)Rq����Z����"������x]��E�Q�?��Q�Zۚv`6`���V��k��I�Rdb|Ԧ+$_�j�3\U��@���#{G"((�]Mb�k����^w�[�Q�%ܛ�>�����d��*�W�u�cD�t&-� �i��(�um���55�ǯ�+Fv�(mD��=8�J>c�:�K�o-��/(���.g 8����[��p������G�_��o!��k��Ma���64l��E&��x���<��^p�e���Z�a��+��@!�8��.c#`z��k�R\�EQ���I���!~t�<��5(9vő|<ӊ<-{+Ti���Tz�Ke�v#JQ^f/Yk$�7��A�u�*}�s�Q�R�X�Ĥkf��o{X��>��}_d��k����:�����wP��U՚ 7�>]��+�k�;Ϫ���G/��1$_(��1��1.�������`�E���Pt��oﴄ�몄�&��I���pԓ<�s�*�~�z�l�{ 9��LK��fh��4�����c�����L�h�5�g��~�p�ʚ�Cs*-����'�˾z/���m��7!�o>�p0\�����9�_��֊įj����o�[hK���Ý^ci~�9��H�2766���tZ�Qt�������d�9L�^�m;ү�9�<c}!��W��n�n�p#Z/��ֆP���័�`B����z�>FF6�mz?dt����W��Ѿ�T�8i���脯�߼4LB�N��*���1JtO�rL�v&�o��D���8�K�g*��KΏ�%��{��Q<SugZ"u6�W�X$�s��C��d.ii��0�����F����7,�v>NWT���\8��sJ?�g����<����iw~`	{�7۰/v�\~xHMa u��bkܶv=L��B*��2��V�'r�U]������/�h8kѩ{L���e�3_�I+�g�1��PVҖq��p�\�L{�b��R�Aš94�4�/�S�%�3��XXd��l�&s�6(_���mk�#�Zƃ��m�RD*,�u����&��d?"L7�䭖�(����>�����B�f�;�q��"��c`�H�9"h!��N�ƫ�e��Yr�f#������͵�c�,c�7?����͇;���Z1�#tm1�qà3�S��PͯwTk"����\�^��<���>L��
�T�r�>��W�2�Ʋ@�A�y���>�����<��Gc�F��1M��$W�r�ԁ���d�� *CMG0�����;�w��'i�v���h����H�g�p٦���
:,x�Ŏr�jj�g8�p��ms��T˖�@�Y�ѳ��eQ@��i`�o�by�0�7��@e�Xb[}�ҹD�����T���.���9r�Z;~W���� ih��Q<�=
����w6t�~���Wց��SL:]"�"���� xIu�BZn�4�,��?�|�t��)�=n���]입�g)0����F�E�����)����#��	~�w������4,����݅
�R�:2��u#����^��=Z��G%�3=�6&3Л��AbLf���l��PʦE�塋#NN~�Ys?�ĺ��9�2�۫E�2�,�'ަb��F�����H���x%x~��MN��}T3�R��|I�H3rb��M��������V�ܦ��P���U'v�k���ƈ�?��Vħ�����x�o�Xh��M����wiZ�������(A��#�*��m�v�"}����^1D�NB��j�כ��"�#?�w�*�K�OS��C�҄?�0,ހ�껴dA��-D3�E��q';��|���x�*^%��[|�u�/֙(2�	GeD���/|�jN~�b�����,x�bn:������{SF��$ȿ���#埙���C}��f�����=�����b��}ӯ����a$�����g�h_	J5�\$�K�Mn�x�3��O[��o�����=5�?(Ɲ����%|�*�'&�7�W��H�V��8�]}�gZ�B�+�*A�=ҨL���>�`˔�`��=ۢ^\%�E@⑓+���Kx��X;(~m�� �|��(iĞ�Ev12D�HH����+��m@�s-��O{�6��߂*V�f�N:���y�RX�X�u3����#ҳ�if1ȥH���k|n��o��޽�c�������C��8�a��H��4����nqa��=��q7�J�L?��J��b��2-�4� 
��A�"�C�@�oꅕ?S�hk9�D�'��2���ÛH���<���K�ŕV��S`�>U���.k�	�Q����"�}Ӎ�����F,��6M�H���-���k��h���i6��T��E�r�P��Tƞ��ń��]a��y�N}�N16�wy�X�f��G�;ɭ���� W��/q����h��dj�իԱܘb�?���H����<�Z�Y����:+��@پ�gx��!(}�F�})![�� 
M�g_��l�g�A|�?�?��m�N�~�m|I���6{Z\�)���E��r;���*��k�!AI½�j,���%`�ML	JOZg��Se���f��ۛ�%�E�>jU͕�%�Me���O0e�����-�2L�&���D��a�79C������|�?G����Ȳ-C�� ��Ln�_'��0v'>�=�rN�e�c9��Ɓ%Vk/�!za9lΰe*�G��4�1>�u�sq�OBc�L�uA���^���j���`�d�����74����.U��TJ����gHJ��x�.n��]��A�&C��P�y���xjƤH=�Bzi�x.W{���K���� [�Wt�Z5�����K}��Q
~r��j�-��K܎�wmؑ3}˦�O���Xr�(�~��;Eİ��%�����9���i��mK���#�`�1��Co������5�nsd����<W}_4�.��Ȕ�'�q�R̢W] ]^#NI2�+��>�94G�E�GS/�.�ZͭQO���Y��x�m��ׯWC�3&)�J����H�h����۵F�xq�K�F�Ie�Zk!��1 `rypo*5D�kb��B����O�5N�|�97P�^����;���a�,M�t��1,8���
��X.H�nqt����c%&�#� 6�h�-���.�T௘(���=�E/�f�*^�
F�`k�\v�:�>)�mښb���?�_V1 ���rи��"X�~ӡ-'����4l�rL�fʌ�=�Z�f�z�jy��;�#���&��e1�U���`���D���®=鵂�h����g�8'���<���H�
�`���Zz�������xb}J�w�����Iٞ䏑@@`6���b8�$��F�&�;����I�rF��������<3�V�����[�H�2���S-��O5~AR��ԭ���.-����s��6���/�A�sy��3�7�s�c��م,D�{;v��ѐ#F1G��]q�zڲ��å�	��I 2���\@�չ�A�j�J�,��&�SH���N�є�r]ke�6
G��:.,�����m;|�4N�����7��gJ�Iw>7��t=s�(�3Ma3y�eێU'ͦ���ٹ�̬ � �ͺs�$[S���$B���\�`��z��,Duu�����g�6�66U}9�@z�ϡ��D?ԳC�t׶s�8�R�A�s��7i���<��v<���R�4�b�b�����[�>�m��j&k��v/9�&{0��gʞ�>k�EQ��,F9����Z�;�<������F���P����Q�����m<����=1��6�h�EX�9[��1��-�t�#&���b��)`:�l���:#tE$^8�O�������۳j�A$��2��&�u�t�U��/���E�X��~�*}j$��6��I��)"�%��2ÿ�J	�hAr�.��'�^a(���5�!o��'�rEl�󩭌�~�0��71��d7�Pj�]J�PKQ�p��%�M�O���暛)/�;jw��C�0a�ܯȖ�Q	1��^L?����s
���ݱZΡ"���œ_{�h�V3�Ļi����}?-.2�������A�aﮫ�$��Sr�F� h��	?;%0�_�C��by�9knM`�T����k+�����{Y%2/	x��#5֮ ����33�� Z�/��i+ͿĻ�ѰZ�s�9aK��������?*�[�r�h��=�|I�#`Ê��{�벏GmB��������]��o	�U������X���j�S���8��w^lbv��*�Qi8�$P�	���\�����-���0�'H����ޟα�fU��Kp=���H�ƽ�������r�?),b;�R�g�����Ȝ�	x�ǩ�1�ļT9(��������VnAK-zx�2f}a�����)ɍ��Ʀ[��1�P�ydUT���T`h�Qm6�+�ӌ=?/42����=N�גl
��h�8�tGχ���8br!��\��C�@�<@�?�*n�v���(P@5�9����ʉps���C�y�<F+J(M����G@���	�6B%q��� ��ܮ���n��#��AUL�ł�'�7���Q���J���ڄH�{���ǘ~U�i;WK�UWaG������5��h�����@paW��큘����п�͙�_w�gʿui��]�6���jTq�g�R�U��L{v�
��������7.��wT<��X�.�5+so)Q��eoR���H��&�J6z����?y~z�B���m�{�z�D�جx�B�^�Cv��2��9�tH�'�!��;��x��|���$�Qs���HRƉ9�J�d�Y�;��5oU� ����8MMx~$�7�o� M�]�s���l�����"�����yި��Rd@����Vc/�<���$�d�F��1`53I�0֯B�hj<��w�ػ�2Ĭ�5�W�wE����Tn�}G�K��書���wF,�r~�����Thꡪ�'���{��@��o<�c��ow(ݽ��Ko�6pr�Wd	�
�>��f������AOKH�3.�si�~MAY's��d�=��sۥs���jq)���Ζ��c	4���R�s�Es�f�M�D� ��0��-�X���)�_{be�"K�$hDN����)V�h���F}�/�j�ef=���C
)��,�!'���p��?}����|B�6�
�3���P���S���/֦��*���5�!���_�}�8-����%2,!EU�d��-���o<�}�U��;�� �楚�<�Hٚ{��G�y���/Պ�x�He��8�zn �W�CVp�E ��?*
9\�؍Vûr�����F�M`�V��a�P�Ȭ���W���se�������Ru����4��7P� �M�%�C'g���Î�d�t�������I3v�����QID�����7n���?3�,�� ��P�ui6�P>����|��G�?�xMkDi�5!�,S�^��ē�����Ի�/��dZ��x�?��;=9�w��ʉ�>���!"1FF�,߽#V�ѭ��	2��֥N���?����Tz��,\���-p0��I��y3����1���R*rY]�0N�!����Hs��ژL��_�s���S� �}��(��`�V�q���Yݏ�3M��?#b�l?+���m©j��{q)F��ݫ��%��ɝ�J�|1���xR�E�;���k�������fb+ї��F8�9�	
b9T�3Amĝ�>����{Eg�_'���~�dץƦR�*��ZX͔|	۶��m �)��s᝭C z)��ޑ9��������rI��[+8ΐ�I�J*������mxﬀ:)A�C����� �k�(��5�u4�8�>�kM��
�+�p](��>
�;�$�0�[��1��S���7��_�j����?����PJ����x:ə���m*&A�����$�6��%���O�i��b��=�6M��ؓ�1�m�Q\~ݔ�kF╯��q�#D����Xn.�w��ɜ�!��P�ݧ�Gg���L���yo[/d=���8�����{�M�-of��
�(�����ʯ�FAB
��yK�m1�����Y��/Gz�i�v���w�Ƥ>��@<��^z=�u�����l���}�s���!m��Y�!������Y쪇���2��4�H�	T�8�|~Ixf9~�-��?�őa�r{�.�`����W���L��O����Fd�>� �_��/��\ʓi��G�G\�P�	�ʋKT
ܔ���dv~�@B�^�JZؿ�8/M���H�ݞ��Ÿ�F�V��/G � g���z�`vLe��ظ�ڭ�t�wE�+ �Q��m2�!�nK>�ʁ��b��_��WFD��9x�ؽ�)(Uk8����%]��j.��_!���4�튘I���V~ZS&�[(�!s8��.}���*8u�n'^��
a�fc���O$�(����*8��GP|Iɕ�J����p{٣�j������C<�:a�li�|t$%�͒������_�b��u���z�����/�L/���bB�C#?Cz�.������̂D��ve�<�!rth,��Ü1�Hb��d��;~7�oߵC3�K�(я���i�Ǜ�֬L�p_��.nW6�|���C���E9�yd�U�-P��dz_�=��᠋�k|U��������G8=� �$�`��z*yK�c�$�c���ػ
��3��B)%W��5��x$-	g����If�ճT��F]c�����,��Ie�C�7���\`�Y�@n���^� �I��/�yc� ���-����pő�1
���b�Ub�����M>�!�)ė�E�� 鶢�xZ�r���D��
�`#B�5��ޝ����pš��MT=�i�D����0��x8�Q���z��,�B�@[��j�>`v�N�:��8�o�����1�Г1;:�����3F</�N'�j�u��=<���'�"��Ki뚀V�xu�[�9w{��3�UX|���k���O�M�|3H��M��% ?4<��{>�_����i�#�gJUE�>+�������/��yK���bg�E����I&
4�y��T�Ҿd� �"�p��7�4�I���i��4�4�"�Kn�.:r��W�N���H^�M�9@�����+ϖ@�֎,궛E*C��W��ϰL��1OҰ�����0�����m���nH������ꊴX?�P������'��>�0;��� jd�ޭj?���⠰�T��ķ��ڡȴb�����~�k$�O��[���2p�o�8�1��u����2��bԧ�@F{�ɏ���'u��Ŭo�Or�g!s5�k�2�u�C�ż�p߆k����])[����g�ɘ&6�yTDoe���r�s���,=�F3�����X�,�yFP��R���R
����=�t�#���ُ�U���:S�*�����k�;���1�9�|�߀1c��d����?ڈ$�Kը��C��*�L�~�,$��ڈ�d����_��`������<m�� ���+�	K���Vh�7��8f�Y>�	1֑I�|��;J ���Jڹ��R>�o�����{�J���k�=޲`^�?B蘳��ӍWm]ӹ��3/�I���)��6��Ŵ�FV�$�Wqr���|8��g)����M�p7�1&�}�J���=�p{��	��,���(�t�
6��ځ�NG�Z��q<X;m4FF��xc�wŎ���ٵ���ȓ�T�<��Y�)͵�oNͽ��w�M�L�m����J���3`:�@VsR1xE��W���{��Wi��V ��P4�	���ZP�ٖ9�˫ОKő���]�T��/grjO���V_��~��v�:~��J�c�`��p���7*aB���H�����?��8^��?D��Q�	>"�ڝ���X�H��bUr�^S�]��`B��(���=�}�*�E℥��ڰڲUZ���ch|k����ό�愊���t/�}��p�7�Z�ܑ��\(�_�)J���!�z�	��	Ii�+�gr���l��D�C����E�'�Dx��c��&����-v밥�N�_!���O�}���*g��G��<M���΂��m���}3��5�ʢ$Y=G�X.���zW�E���W��b�.�$��B�Y4P.�m����j���	y.�c��mM����IS����K!� D�{�M��M�d�D�=��N�&�L�j��*N�|��Q�v��!m}K����!CfS�K�k�dP`�a�a�e�JT��q����ux�1�/}��@���1*�3e�lJ{~�?�@ۨ�R嬧��F��LAC�gg��d�zMd��a/��}!�1"�a��
H��h����)8ՈW�1��W��Fߍ
9����~��_~e'7���)��h��n���TFmjE��������(P��]��;���9뢑?�qP>��d���h4U��i2'V+!y,��z�����H�Ҳ��2����,�!�c��r�_�cVܽ�:�G����v�F����\D !�d�X�w>��<�����N5wώ� �N��o��#��c��Aؒ�s�K�*��\zS���S|�{�NT��+N�u�)��ľR�ze�S�@f�Ώ��j���c�w|�6C���H3O ��x����$���m�֥�m�KYk�^�����[ڥ/B_k@g�FG2����x�8�����l�Dt���c:�-?Sſ�y��x"��4��l*��S�t+I�t�4��?���Ε~��H��4ƚ�q��ײ���?1���\O5a�;O3cf�kU�'w�/[�'�	*]'�f��������KBx��Z ������,^H�
QeԒ��M��\1�ΟWX����\uY�W�f��,*Yn���T_ۍ�l�^�WG��6���2��[	!`-_�O�� ��,UR�	Z3{J�g��DJ
|DA�^x��vL&�����z-�b"׃��>*�1�0�y��	�cq��\N�C���\	@�:AP'n�Ajh�F���YN��%l׿�?�b�����w��`��X��g(|���»Ms�VH�e����mK�&fyKUǝ.c���$晽_��4Ҽ��Л�X�e��M5pL��` �7�u��R��y���";V���r�o9|j����A˖��GK�s#�liٌg��NȺ�o���K+��[�~�1A����t�X-B����/-vBzĻhQOB���J?����O��O~V�֟|����C�HdP��y�о�O�"�������م:�k�����.�nK^���:s���A ;��(��c�Β�/�O�41�jj#B�z�-����V���c��ԍ��r]�I����\|����1�����w�sy�ڃ��N����+H:D�~a�{7��^�B����e�-�Q�����RWrc(
o��T���Ut�ݢ�VpN�jv��S�MP__@	p����-f|#���|�.$x1-N�'1�Ma�!V��x���lKsSu��'�>�m�pμOͿG�N�M�({�돋��a'�Fh0��+��<]��Au4ʘb��J���fm�n=��9)��Y���{ZtP���5��/$�����i�M�"5���>�{T�n)�i����yU�G�I�\��?d!\߷P[���G�ﷳ���G5��=���KG>�<������E�y%P�\�枻2�#��Ea���6)�T&N�#�K^Hijz��%P�$f���]~l�{*�g�?BF��?UG��Of.:�����b�k����T$u���6(�3�+.R.������*=�<��5m]h�X�0���1�s�.�s-�5�����OIP��&�j�j9x,�m9g�C�&Q5B&J�ҷ����Ě��
.{�dL�N��AC�]�qF9H�E�ehe�� -+rT���Ҳ`-�	&7'�����npI���?+�k�34L��s iK�Tn9Ar�TI.���EC|0A��Z���7"�L��Y�Y����6�ڼ��t7�t�⠹�:N��>���MX����_�#����?nFë�s͊�����C~\���� .ɿڷ�Vr�aH��"ɛ<�K���n��Na�V��/����%�'I�}.�[��!��2 ��`�\ޢ�5\޷�B0F��]�*�2n�՟e	e�'6�/{�Ͷke����S-��H��>�t^�"�E��
�p!����(�8^*xJ�����+�3K��)�p��-+7&38)Iⲫ�w=yn������ �@�f��}ʻ�A��S����"�WVHL>|���&0��P���%�~����ʑ1@�J���m� ��[Žf�a�m��A%���q����+Rp����1�@e�V�Jg�hR�_�w��6��O������ۻ���gTx������c�?�X.����� ���(c����X�����7�˹X*�ꄋ��.����֭����o�[��Q���`$�a�U�Ȼ��>��\	|;�v��@Uŝ&�و����?�a�!\k�r�W�l�z���g�����rq����K�����ָ��n��S������W���.��le���ۼ��
��#����
�8TS6�#�0��	���ע  ���*K��B'��m8��G�e�E��0�y]�	��:h���,-�x�k��Z�T����NTB�dU�Y��k@đ�a�)�O)㸚��r�r�FUOV�Ќ�lA�u���j|����L�_ܞϞ�D��Do��6�7+?�`�AkUw�O�&�ۇ��i�hR	JghA�~��ۢ�:�Z�ف���ޚn���q����ٳ%F$�Q=܏�4O��9�L�0�1�N�'�ʣ���j���G���c�F�P�>�����\�w�?�7����1�I�L�9�";2�����w��C���T��Zӎ&����[[b��v�GdIsg�
�������sm	��k��x��F�r�FC�#��* Se��-f��m��E'��<a����B�����H\I`}��S�s�B�9~�Z�U��v��I�n�+*�)�S��{d��}BWd��2���j�������	r��X�F� O>�l�-!0��*?�m{�k���ǅ9R�'8�^X��ӡrW���5F� �� UB�vA��k��	�C:�Z{;?b\�}�Z;$�|�.b6?�-\գ�t�s<��tW��ƶ��J��O��)�XN�Ѹ�����s'�	��#Z��S݉m]������W�7j��`�������v��GK����bZ���pCf��"i����F@���赐���#�:�1˿*`���]�&I/�Z�c��֗������JI9	扤&��R�����'B�ѹZt�*�V4W�\��͟���Z�	��H��U��b�y���Vr)J�,�?%�U���P�H���҆��V�����=r�v�L�$$}1f+h�����X�pR=uj��]�Z�@�����>>`ۡ"��,'�;��A�Q�P�f]�!ñ��<1����p�H��]�.�Sk�I1/b�(����r~Ԡ9gi�q���X�b�|��ߩ�2c�5�cO'����Q�k��hΣ�vٹ9����?F��UON���h�C�-�ӫ���EV���G�f�{i�*<F�>�b2�tTl��!S��.�绡�:�N�pH���?`�?)�6F:R����4��%�Hk�_g�������-�1�����#@���誯�I�u�*����T�<G�x8f��M$}�D���E(y9%��90_�E��󉦭T�P�(���X��s����n0�j�.Qߓл˯g�V�����'���tՄN���>?��:���\�M)�7�w���s�ש\� q�Ɯ��{��_׏aE�Q�M�	�8��s�1x�vh��iB�2Zc�'��9�Y[]��N��%�F�������s��կ�i���	C���a����#:ŠH:���C/�s���~�{��R�ۏ���}�E������϶�rR�^��B\,;��wH۷8��jN��������?�e��m�v�}NC��O�\�N���H@p�R��Qi�5�7�5�?��oYY@KBp/Ԓ)QSl�(�������-�����\���^�/���9u�a��#�Q�I���I�p���
+/�Lm*ϡ�76�߈�q�Xr�Ѹ����0�ʹZG���p�������"�a�9�s�&��8 �vIK+L@T�B����$�t�����3GgD�p�$Cpwb_9z6B�v����g��c������\|Ӓ���xs�$W�"��K���cr قuܠ9+��Ǹ���
�+�B���n���\7���ԋ'�T`�r���Q�
�տ­��I��� ��w$����9,^Ӯ�I��1�z�0|�5����a�-|�)����e�: ��Ǒ���Dqʎ��Sѩ��%�M��QKE5��L��<�aF��x0�M!��lya:���%�S�B��G>J%
�b�؛�@1�;0|�}�B{�B�Z.9�9�2�B����SN��2�:QO�����
d$���C:���E�<��J^xF�>H!�n��&�W)F.n1�+�r�g��M�j��
>&K�s�& 2��ce{l����ӻ���c���v^��σ���6t��c9p��2�S��7�	��%��9��@��Jc���a��S|��C�܂�/������?��O�����i�1i�w�E�ziK�� �8��o���D�n��$�A��菺�ܰ����	�X>t�#b:�D��+�p3��&6�V7n�xN�<[ݧ����ZF�v��Bc����� v7b-=(�`&�c�;�� �:���P��3�������d?��Odd�.Br8 �՗Y�i\&�5�P�o�����*U/��Ndu[�F|���Z������Q�fN�l��ߎ�v�P�V�6�d���wA=p^�{+4�ׇy� �'g���M+��G]ofǑ��������"$x��X�^3�ѫ)x����$ƙ�R�ۖ�d�a��?7"�@�ٝ���3Ca	��4sX_�?��;�g�7�a��%{�	-R
��ׂ��H�3+�Z#����T�	�aA����\K��<g�S��>X���y�lЛF�&3��m�?7G��B�K��`D�������G�|NeF�W��;��WDrK��_&�Q�ǣ�`*�kA۰��m�Ｒy>+���4���̂NA�zg!�ɛ��s�>�v�8J�Į��1.$�j��o�9����K<���<࢞�I�&��9C�Gm���6G���Cv�uK�m�x���A����*���e������}&cHn;�pт��x7Ш^EVW�n⏙���Q劾�1?��}�ߤ�a1�(��fx�BXMeM%6�NY����Õ�#��y��^Gck>i
��:�`��S�qxcۈv�mrk���Rrڟ�*l�m���#��x�X�\���^`&4��p�p���e�ρg2�p.=�]w 81x�@ca��p�F�Ps��0ڰ�Ujbv�{�CF�u5�L(�`t,4�j9��U�'i���yS'�^r�
YS����.p�a�+�S���j4x���j�2B�M�\ �, Tgx��b^��61�hהuŋ=���Ԡt;n����e	�Z�)��K������K}�B�������	�2�������8ʢ�J��гd���oB�A�K�`���h�'W��`��ݻ�|�nޓ�g}�p�D>2P�7�m]�k" \E�u��v����"�e`U
$6�=v��	��W���BQk�4������i�1_���R�	�7I�� ��`�#�f������jW���n��\,|��
���T��
��a�5��'��A*nsI�kg�O�y&dSAj�~��bC����+�.;�v��^��D_���5"ĕˌ�}��a�6��(CEo��%�e����?��	z�H
�Q�h9����إ�zVBȫ�� �7�Y�+�jK����>$!=$DN�IXu���M:4��mQ?Q~T���@j�x�3�M�o��X�amfEX��S����A�˻G��}�W:�.x�)Xr��2�z|`_T�������ŽQ������T��m�G?$��g0��3���
S�<B��ͦ�[��L��}��Y-�rU2.���y_���@�iۍ�P �N���X��Kl�l�٣�̀�iۃT����T|���8�?�t;�r�	z����k����iM�z�����3�R��;O���� ��dϿD�=mgRI�
="��}��˹l���2��%�}�i	YÍP��Z��/Lb�!xN�oͱ��ήP����q�L^z�.���5h*�mU�Hc��t5['=����y��&��K��j������P�^\�#kM)=��h+�Q�.�0����Oa�L�y%���S	aF��!uBD��a����!?�Z$3v��� x��-�-}�0�,�tg�L=�Y�'��$޴}�,8{1sa����&��5��Kl���(��5�r�ϔ�?��Gb�LZ
f�Vn|�)D���ȶN��
/~�X�o�ݛH�.��+�6����Ç⦳��K�l0?;X��D���
ɦ��˧ʨ�J�f��/�~²�U��J3G�<�$��\A&J�/2����̗?���h�\���P�R��@����)ϖR�����ćo��
�ū�=/��%\f;D�P��V*�9������b��E�4 zVp�p>\�nP2BW�%C�U�D�J���ɾ�"���ۃ9����DK;�X;�p�%��}>C��n��1%jH�q5�X��W�`�ħ2��)�Eb��	�m�­�tɭ�yˤ��P�Mc*Z��
��	*�010M�d�o�CnQ�W간��s }Ws��GIV-[L�!���q���.���j��)H��'[��z���û�Y5M��
y�@�U��)�}��L�VDg m�2Q����{��U� KG� �rξǀZ���LM��;��O��)�:Q60��|H�M�)���/��g�qwӟ�&��?o�c�����*Ќ��J�GR�*��_[�Ս=x�T�"
Ѯ7(Y���
 ��&8.z�1tU'r���_��;�
��*t�Ge�c�jV^��pj)z�A�\����@a�er�NLAc�ގ��o��7� l�Д��&N&�3�4"W�G��X}]*3��B-֭����t^�R��6����-�Br���xz�����hӖC?l�=�,Z�L����Bэ�~d��l/�~b�}T#d�Ǘ^����-/��s�Q{<�)!�X�S��փeۚ��7#.�u�|"s�.k���P�З�i5uu.mI)0ϵ�%6a�rr:��&�zA�[����Sl2��V�����a����BnrG�y�7��a��z�ƴE��96k�5��q�;�Q�'"B��O�H����ߧ�J�$���,��9�rԚ[�� B��t�|�����.AS&p�2��+! �����⪹�6T�_'d����M��d�x���w��AvЁ��SRt�v����ަ��Sa�� LU�p�#M���òV�`�w�<��bq� i�7�j5���� V���
����F�ml��$�a��H����uhY�lW�'����m �?��\!���~pm4��_d��E#p/'�>�ߍ��-1��Xs�ri���G����p�m�5���ɵ��W?��2u���OX|j2$[�敳�$�5�ױt��W#��(�O;�7?N�2	�3�ڴ�G-f����뼔T�S-ϲş"k+��9�C`��+�o�kx#��9=�������׃g��-A�#6s��L�Č0�/)w�Ҭ!�j�.��ǲ��T7[�!�]�+����_cWS?{e�Nm�����tiԵBj����jI�ɥ%�3�XkE�6�UȃOj�Pl���E2t@��T��x�A�gHuߏI4���ٻd�����"?7�f�d�~��ض��7ۑ1�x@��Ix#�~��	��:x�oĒ�t�P�Jz���G;�i^hO�G���m�VR�	��F^��� !+����+��ަ��)Ncۀ@��>u�軞���=����Эն]c�7�x��@��~��)y�7.$E�e�F���Gա�zг[�B����$�sTWT�'���y�	��nv�(�]=�Vb�~�׮�n���B$�ד[6r�X.�'b��53�e8u9�i����X��p�4�dQ[\�p?К����,�֐��{�;�f�c�_Y�Ų������;o�����]���B����g�:���^��OV9J9x��lr)'SG�Xe���:Hp�Á[Cj~�}_�Rm�+�ę������� ���5qlr�}�f��8�+�75�6�!U�H��ל+�n(5�f���X��dV��3>LE1 �哃҂hOi�JT�*��nN������M���ym��#��G9�_��(-P҆H3�W�V|,�%܃�`��r� $C���%�Ϩ�=s5�4KB$F��B�R���ڬ����tD��c���/��������"�svY�$s>���U�.�(��^�C/��jx�����#�8�I���sc���y9b"K�&Drݟ�3��}̐B_]H���̃}	Q��^Πb|�U�Ј���|u`Bc�ɓ��]���18R��
�$5�Dx��.j}�H���E��8��`qo����7�-eey�a�����í����؀s��sKfp�qx��n��A���?��m�GT�@Iwƙt:R���W	�*n�&Xq\��L���T%�S*�)�&nF
���Va��Pv�T8�9&=R���(7L�h���o�!�K�^��ԍ<=P��lZk�R':v�e�l��+H��QΥ��<�^`;c7����sG�o���)f�M��F���3��l��8�_�QB�2����6c�2ܴiW���5�o��(��T	1�ԗ5r:5�B�#^���-�0�?��v�#�W5����nc�:�H�r���P�� ��9���֢y��=�H\4�>ݎB��IH���3=�8{XF����Tփ6Ӡ �R��0�����{u=昡�Q��CW �?T��zB��]TI�rfm(o�B�s�2}��T��<rxm`0Q�/G����,�^��U�as�� ��vO�A�ޙ�9��8!�p�����'IU��w�[?��5\���幏�d��لMXZ�^�ɍ����Wt`���n23l���-a��$�̎Vo���Aħdq�҇&_��{ �M���	�.xU�f�<���Ĳ"��� ��a�+=�\fT�"��v.���*�=7�l�v�6�\���..��Q��:[��r˱%�OS��\�֏��*s��NYd�=�0��j�a�%\�U�NWf��<�A�Ο�������Y��������G0�8�}A�(F�i�C6� ��nNBj�h�s!�T���`|8��d .��Qg@�����n:�)���eW�b�P���B[�M|��Ky������#H�q��p���D�.�1$5_��O�~r��p,�
&�U;p���Raҳ5���z�o�y�E�����	��Ɍ)��)O���d�ى�O����_|���h (�Y,>|:��"2��l�$D�饡;�%�e�(F ��1���B:�#}bpd�!�
ά
/�C��|���"�
PT�jx�J�#%�����J=r��;���\w�C���F�*���9�Bq6�@.�2�����b�)=b���Ŗ�Ն�("���,�o���E��,��6�/C�V��X��0ct���6�I�c>������j��|  �ܵ|~»CPI�4M���kYeo3.g:#y�_�����A&���;e��CB�r�,W4y(�B�
i-7����F���{Ӆƿ���A�7�Uu��S��Њ��o�:�".��z��=��D��u�ܤ�o��)�?r%���6�
�켌C��IR�T���iAE�ط�n?�ت8^Q�B���XEґ\>;�A�J$!��T��Y��@mf��oKAm6�O�+���fL�	�Y� Q�ɱ��Kmf_U�j3����Ԙ��F֌ҽ���������Y�ƕ�������r�h'�J�A޶ʲ�YH9�a9A��EkZy�C �ȆT�nEn]�:��i��m��ʻ�=W*�]��G�KE*Ɖ�R�Zw�����p4���8.�#����W���5��)>�6��;#��)k�l�c�$+.��GrWU5�S�MzYa��iW,�ǀ��#G�d�;L�\P���5��!��H�=����`x'5�#�f�R�w�'eP���1�i11�������:��cר��^�HA.�-���/)@5-n�k�T=�j_�"�p]��T�No�������BVf����H0������;�p�lۮlp�{Y����̪p'��(�q��-G@92E�l�W���������VU������f
6�1�,e�0��b@o�.C��tf�ei=U��Eƾ���q�rp|��°f�R)��o�,��9����9;Ά}�i�!wO�H}�<���{<d��:�����'��(���gJ?D2@p���ܾv�{M׉�?��Q����?�8����$+��F	i�&�Ml>͡���=O�}獿,Rqu��0��?�d!�D0@W����U��	Lt�
!B��lO�瓾��^�g�ն�V�Bv�mG�J�N��]!��9�-m��?}��i�/�Z���һ&���&n�f7X�b��9�oB,�o�%?`>�(U%�p&A>M�n��v?�$��,��5��OɅ�Ar]��3��A�č�MZe`?&�2�b�7�g���~�H�|̖�p"���ܤ�?���:�|S�<?6>p6'��+�m�8�x'h~��	�C�?�4�rE�t~2��-�N��/�4�ۯٓ�CZ8@$�7�4;#�sfɩ^(�+�r�E����<S�T�e�lx�#��9�ARǨ��R�@�0��~5)w� ޠY��J�*������?޼2�6���D�t�z�=������`v<�>������΄B�m;=Us`'�x��o� C���~���� ��o[5ޒΥ��͖2�Fp0:Ki��miY2_D�(~<�:w
�N*��5�!��J�B���M�T�;�WUFN��r���L������Q�F���ݱ��N5�$�:QsΔ�Io�[�>�)���'����%�C` ��-T}����(�Ri���Y�K��m1��o��h�LY�O�����{U�g�4� �XOp˗��|=*������W��gs���S
tt��?R���,ທ3mf:ؖ+���ڪlMy��6��j|��d�kO	X��T�
�ҵU�㣠�a�)�E�K0�D��4	Ĩ%z�C��j)�
�\��!y>+���~��)Rn������1u�����'��<�B��.6�$�X%����یfYg�5���Pb�����,Y.��(����w9B����ʮ�TE���Z&�G�$|�-=�I#�?�Cq�v�^�d��AQ3@�30{"� �	�z{����˭QV�Q��O.-v[�ڡ�(A�X��e��ѱ ��������/�yi�Z�QC�&�|5����iL��P&���8=x�2�����EP��S�-�4������I�	�bDF�Fz1�� ��ÿeWh2+f�C�����������o)K���U�E��_`ɽ:��3"��3t�x�in����PC��7Ko��*'���<����7*'1�p���̿CQ��Lڊ#N�1C-��r&s�����|���B�Q�뻷^<7��Ņ�S��"N�Wm�n�B�Rg�\8�a� T���v��n�U$7�P	�4+�a\�Ma;-������LX�񎷚�k�.�]��S�g5��,m���ʉ�}��"DH��R*��<
�,(�{��?}os�����K�?���VQu;!����D�����5��Mt���a^6��Z����ç��Nx�)��F�]>�x�%�T��tð��@���R=n���0W�`4]���-j�<n1z��@BpqxG��O����<~ɟ����?��zH�.%�zS���Ԑ@ߥ2��b�Й�ڟ�9H� �)98h�92c�T�5Mcv�>è�t[��޲;`e���(FoD����e��fIKS�x82*��I��6�0�8�Yf��I(a`����oK���M��>�K�z�$N�q����&���X���e��uhӦ�և�9`�x�Z,���:��X.,ߖWo]X�xA��~J&�
Y�P�f:�V�{H�c���x�Ս|l��a�'���?[ViqG��%bV��dK��uv���/ۦ�p
A�B���@�CxH��˕�?�m�Gg!���T�.�C������,��d��]�M��&�l
/��9������]���!?8ʛ{x���A�d�{ц�c����DW�75�pj�LF����#(�%��\�@k�s��JE)����^q�> GW���>~���OI}��1PӰݗy˙�����i�qx��UNU��o�[Y�)0ȃ�/	�����n�%'��S��~�2c�j~�)ݥ1NվxW�`��qw��oъ<��j��]۪��w�� #?�6e*�uDp%%�8�,ܭML\-[yI��fw�����WI
0%�~��U��0�r ���݇�ׁ�^�D��N���x���9ƲE�8A9�J��e.X�]{i{#�,������h��n�Np'�n�L�H�������F��)k��y���wCA��R�*D�W��Ԭx_6�~y+���\.$9����f�
5D5N��cͣy@̈́��쁩.�^K�F����}��e*�'پi'M��׽� Xa�s��*d�\d��L�tt��H�$�{ط�۲�+�%"Q����͇�(v����ڏ���L�y<
��M�Z(3-��<�<1����_��Z�2y��a�5[ܛ�5�MI��"�_�S0	��1:q'w>*ز�_W猕y��$����k��z��l���qygsE�ǔ"z[I���J�b�����uo*h��J�����}S�Ҟ9Fh��w���>^�8�ꁳ�������0T�����	,P3!��j�#	�Vl�*d��gM�M�]*eVU�BJ{��}O���q\4�"�L`������z%&"m��y�+���r�7[h��N� �wl1@�{�DۂN���S�*ե��r�pԻ�0��1�s��� j.���0M�2#�ƍ�����}[3|��N��I�S� ?E!@�uS�+���M%x��ϡ�ru!��e*ҕ���_�!C�Z�i广(��7+7EUj�u�6/\>Ф۸����ɡT��+
�A��N���q���H#����A�����͡�9=�\��F��<�<�����?a��$��\���^X&g���؛S��L9#yI�PT���g���p�f!sՋa�nL����nc���s2�Q;+AԐ�K�c�ݻz�u����D�;�����k]�z ��3^R$d�J]
h���)�h�{�xK�§ج-+�Lʁ?��y{T ���ѱ���@-�d�S�-Ϳy��{�	�;k���|ob��5"�;|1�Y�7�	fz9\���
75j柳??��y��ۏ�BU�f�ק-�O���旸�f*|���|:y?��^C�Jq�=��#6�I��񠝥	��taB�4��x���kƗîH��ݻ��yZ��C�E��T�o��NU�X�s����eŁ� �.����|�� \�H��c!�GvG��6H��Ę4�j�)����	�V7�%�Y�I�Z��ޘK����� O�aBbjb��kEH��4���%\�Ŕn'6�{`A�F����/��{�{9��;táLO+�c:��uk��;��1��HR�l�� ����ж��P�4gՁ=8{��F	AC���_�tWV��ˊqW�1z�Dcś	 7�u ��jM_���"�u����?���c�����*/�}H�Xwڕw	o/�ل�(��)�{C��w����Уp���ܫe��F
<c��-�����.�����g�)0X7y�:��s�amJ���'��x�JpE���J%S7�\� 9�-����X�(.�%��DE3��������aȓ]T����ړ�v�m��~��@A�g���w���,���t�\�<ע�����T��/�_����j��]g�e	������OU�u�=�oI�aˡd㔼�O*>�6�"�gUR�i#��PF���1����Z�J��y8�%� ��̛5�|��*+<H&0�ؿ��\}M��d@qC�ۓt�Ho��$�R����	?�!��
 c�m��@��<H�Rå�{Рթ�А1����Ȝ�O�{i��3�*����ƀ�/�H����*���}QΚ�2��:���.�J-Faf�'ٗ6�w#���� ����*��n$֞�s� ʤ�G϶^����r�5Cup@7�t����P��?�isWJ�9S�>y��C1mN��Î�+�+�h@���v�`�ô���k�hCE�*���Y�>�o�P�����=��ΠH���&o,�|�nN�7��8pfh�?R���CI���x$�?�&�3�x��z�؉9A�U
h_���Rwhc������$���{�>��pb��`Ze���"���
D�bC��c�N�Uǔ%݁W{�Q���x2��|+��N(k��)�_�,g����cXt�>x�!0
g;3�1.8�O�鯕�C�<'�H������L{�����#5"aXܤ�"-�,�p����C�"�V�%Z�]��d0��i�7��m�����`,�|}�˝8��E�
��y��)�I&۽�C{�=�Z ?��G/��f��VIj*��Q}��=�p�r�����<�U�{���=>y����rz��ϗ/\.��JAB�^��c��6%i5¶G1Q%�����w���,ي��̷몪*W�<�M�U}�9�Iؼ� ���z׹�y�����/S����_V�k������^#�lU{�cM�C�����?�>g��HC�IO��D��],�A�vӤ���Q��Q�i����G�z\���<�O��ipT�� �^��{bZew�X@�����Ϡ���J
�t'P�2�3R��me�8��� d +�YS�
��e�	��v͑uM�N6�ܨyi�31��g�2�+͜�͈dd��z8���B}W��[$�����``��G���=O�W��F����1	�����$��Gb=`�.�MB�c��\����7��,�	~}x��wK�c��soe��̽U���cS�6^��.�{�d6��Ub�f���?��z�45���ϊJ����<�,�b��v���u�qfT�E?&����0۬�/H���r��Yh߬�F�Q���:��oB�ʥ�N�:�DB�F�hIaWO����A}6��Ҟ�w���K�HyW;��Ae��b�5���QXC%7�dXg�g^�Y�ɩ�u�8�3D���.t��G�ڦ<�Ẽ�Ջ�Yds�//F�˛H�qF`S
0f�.��zL|�\dގ:�����/^l�&���a�Hq4_�ZF1�[gB�.I	��e'`�Nཬ5=�@7I뼢j+��)�:=f�z?��#�� � �rA���M�",ћw]2;��í�4�p��lz���K�`�X��Oh�[��#ii�ytS_�$����e�J�iElZЙ��8�� �"@:�_�	�g?Q����U2��	s�tW�(@��'�D�7�3(�J�۾�2U�����|�0 ����o��b���?�(r�M���lH2�(	aN*k"��S��3���ܵ�7�C�Z��Z�Z��h�fҤ��+U�T�=c��r���������&ouT�#��%�Ͽ�F���.�_�]��ܯ�ٗ�	D�<�!���2�=�.�&�DD���{�P��T���T�ن3R�L;��r|a�y�~������5ͮ�~
�'F�5��T��m�L5Md��棪���,�?m��P�p�hۀ�Amob&0�(��9ߧ��j���B\RqNo�U�ه��>u	1'���b���Y�]�c|'���x=��f�pDK�g\�h��_9��Ia�I��[&�Mx��i �
�M�T���`P=T�ã]��rT���P.:�K�!�
��@�z)�^�iXs
U����aGz��K��S�N�O#7�����y�	��־�NE,y5��,Zk��"X6�E3��*�	y�S۹�:>�m�g=S��5��9	�kp�4��s��,�ʔmw�/�O��"/�{W������˦�Ԏ2�m���F�WZ�9�����Qݘ�9�f\�&}Am�c �H�-����N��l#��vcR�1�a����(X��h�篅�0��\�|����	��Hu��	D���tn
�3rKA�4E�^�.}2�-�l��~,�n���t��F����l����ք���8ɰ< ݞ���n��>��B~�q>0k��qӄ�a�1��z��J4�~��	ޏ�k�ϲ�R�B����U1�)J�L��w^�m)o	�*"�;�ω����i����/t�^ػў�h��ƫ�O�s��#t����徰Q�p����枙&1B *g
R�sT�v/�:v
����2A1."1Ɣ�[��羲��W��z��iB�Z3{�ux~{g�g,��W�7~ێ��*J�`{�^.[�z�$�߫04j �*�{Ha&2z(I�5'ԟ�\6s���%$=�F3�Q��"���#F�HH�R��TS��� ���D�~�AM&XB?@�����2�H=���H�2㖿w�-�N013,ۏ�6b!���[�Z�
���>����=�چb�_��K;l6e�6���Xun�͑CdO��8��.�?}�|H��qyY���#�ș~ȂE��Yp ��������E��s�3Ma�C�-!�˅�CKv�)��$�����P����F?��k�W�.�9�� �˲|��޻1�Nd��M,@����ʹ3F��J:	N����ao`�,|k ��Z�fO_ %�aP��/H�`Jm?�`�kq��C1 ��'��y�����rp�B+��JQu��-��_�I��s�yN��*K)^��n}�%��r5�* �"���nV2�6�:�3��}��g�5QX��1�n��z���b���ͨf֤P�-�`��YH2:����5A�j,eI��2m����� 1��DϿ�:�\����W���亪p�R�i�ܢ�d8�x�+�!x��X��Ȃ
W������j�F�C�Nß�r�`�^s^ew�pO9��5�d��wl�=P��6׾7&o-+��������m&T�(��."z����	b�1AgP�A�E�N�	BH�Y�M�ݕoH6XM�eh谱0��f�o��� o���\6�.�Ӗ='��'��f���1�MX���I�	�)�H�l��p��*�����Ⓑa;�hB�
�4X�IW�&.%�{?L`6
z?�$7�R&�Ħ4�;��h��3P#K���~�Xɀ.��8�e�r-�����f�(a㨶'J������t��vn鯪,��̊��p���ТE�E�U����~��"�I����S/��ȸ�����K�M�}-$ �a��\=Y��0��=^�򭐲|�q{���.�B/b ��۔�V���f�M#1uFQ�XY�="v �d� �e�uמ���� ��C���j_}�\�]#��d/��xܢ�+�n���꡺>)��.Fm�ɺ�e�B��);���������6��z`b��x�S��	-ٰ�Ar��[s���S�xr�J��`Q��8�n���U�q��@6E��-��2�m{tc���i�H�e"���έ+J� ����'E��RJڙ��3r�`����c��߱h����]d�n����/k)A�\W��Ʊ=�9������g�#�/|K]��8CU!rnq<�`G����l;�Fx���-H����UO$�0t3<����O��W;����DF3��Q	�[lԒ����U�ޝ�^8�Y�T�A�y��t���K($ᯬ��648�##�
^���F���yN��j���ts���T�0_�%i�Ķn�G���X�XR����5�@�!���v4-X]�
3���|h�\�v7G��*�ݞ�d��<���U��T0���-"�,�S1�H"b+�0M���~����ۏQ���f��_E/ѓ��ݚh�c��&� Y?�2#�T�my��{� �o�+�n��BF�a�?Hߟ'�u��ݤ�,�C��%p�qA�$�]�|�>ꐝ,讁��S5��rN�R?4SE��H��N���u5����,ۭZf(����T��L2����s��eJ�]�>�ZYF��_G�5��	�h<��K8㓞��5�∞���9@����bc�%O��Jmc7*��Ko�3U�i6	��:BVvI�7/
[u�tJ%�@f�,#-��'��4{�(O��H%4�
��_��P��/=�Y��{x��P�U5�����C���b�nR�˰=���>�?}�r���N���:y��w�p@f"f�r%�J���һ��+[p��U��$��!���;�jaCq��n%^8��7�~c6���b�O�J�s<�WyI����%msO�&���׹9�z]�w]�Y㌡U���g�i;�=����6�I�����\x4�w�od)0v�$Sǧ��ޛ����x��+/#3u^��6Ua
N�
.��t�4�B�Ƚo��]���Ֆ����9�瞋�]�Gs̖V�n,���b��.JA7/} pi�,c���3�U�7-j/#��bm�`H<��v�LH���q��|k�{>��9�=�	�%;��n�e�}���l0�����DZB�ŌAK3�kR�>�4��g���_]��4�C,����ixMJ&���� �Ľ�?��j�!�3�矄شAe�����2f�ꗾ��X�C ���@��t�,�L����%��,�o�A>����`�q��0Fp&%آ��}�lյ�$I�����E�zC�`�b軴E�N��`y�B�~���`ɐ�s�)ao�ug���~�3+/�~�	5�&�%a���h�{pW��I�O/zR��v2�kM��R�_�r�<[����F�	S�-���b�W(a��YZ��f�x[��? K�W���hTCe|�?M>��$�;O�;�1�0c"��0r{�(� �J�1\���k^��@Bj�R�>3(RN:c��r$G��� ݬ�.+����9>g���������W
'%���ٙ�������9�:�/"�Hs�çaM^6��/�ܓ���
,�K���0����WP1UX����_�J���h�I���=��xֺtƶt�b�ہ�h��3Ьj<�:%˿��o�.=�{���hI�F�� WuY��F��d��T��M5���F��sry���t�x�TvU�Q�LaZ'��Y�Kf�I�K7q���z0�'����.�#'ge�x �ꊁ���!�Q5��|Y�}>����O;�~��7���J֠ke�gc���Y3�dm��]�R�z�q!�W`�7z!]�٢W+���F%i�r����7�b��'��-�.^��e �`�4��W&6��-����Qè�1��ϭ�����7>�A��9q�Hڤm/E^%v��L%#aZ+3�(�#���B��we�lFXـ|D>��q��x�������ވf���:�\VD2��[é+�d�����H]��4ُ��a'��[TV���!C]�s��Λ�#f��F�����8�<A�Z|�]6r���;��9x�z�x��h'������Hu:��smn@8�P��3u�L�mo���<����y k#o��`��" �)�M�/��'���CD9�cs��Z�P!\�m�s$�r"��`��^���˰Ȱ��|�=����d����NF�43o���0� j�AI��� �|!f��;�J]�x������W!]���M�RY���vZ5(��o5� J˖P�-U�,�O�Y�������Z� kk��)�v&�}%b��'
{�1ޘ}����[����e�����_ZW��?�̹�/cO*�����_���D3�W%,�%\3�/+:x
����ט�V5�)��r�6(ʷ��#�[ =��03����.�_��tܹ�m��7P�>"f�AD�0$ˠ����y�]�(f���kg��d;!@�=�ڤ,�n��!Gn�Ӊ�{�/�>�K[z/gŚ������÷�A��1��I����L���8H�P��&�tP��qF��f^�pҠY<X��}��&O��@ңu��y���԰��u��C�Vp�R���l�.�� <�z�N���fm(�9�P@cqq+��4��i��q�rl�� 9�����~�خ��7����-�!�:�C�&d�e��r�mq��7�	��'�y�m���D�qwCR�;|�`FG@�<\>��4X��������� _*��iV.�N�����"x�!@!.p�m�#�(Ӳ����<�G�q�#�HS���E��I�4\��"gX
�e���!���A�m��/��_��k���.��h.�g�f�\}����֜��m�udJ��<���'������ՙ��z=���)�*6�A�N|�^�GT���t�q̪eY/�n�"�F���9{�]
!_Yl�h1(��F<�J��v*~`���t��~|��I�&�����F����6y\��NN��^^Bݚc��hc#"��sݒ�f^�):4�_��T�'3L�3��% 4��`���&u�o�~�[�K���������]��a���[�Ew�+�O�2��ff�M��C:T�Q���(�?3G�]P�hB�&(g��� LH�����g4�]��q{Ibm�ʻ�4m <��+鼦=�mj�s��{��|M�(s�Kbξ��bq1P\s-g;���hg-|�XV�A���:���Zz�	�ɐL�^��Y�!�Iy��M�]	�	(�}k�9�#_��}[q���|{G���kƩG��G�?o%��=���"�}�����p4�a~#�Fu���l��]�El?Ax��������&�(�S�7�eȠ���=~�z7*|M��~��۸R�'�������"�s��VqK���9�_��49�r�p���Q��F�n�R ���z��:��I��q���܀f�Q�c�]0k:\�~v�,�|D�}Kצ���#Ļ��� ��]�܉"kO���8�'����t�v9�������`�9��i`�a��p7w{9�Œ)��!r\��c57ŘƖL�_֥���V ����p��@�C7lE6�C�mƍ��?L��X?.��`"D����	�cR8�1�}��׻,£�SX�3U���Y斐�$R'�4��׷��?p�Nȷ�Hx_�J�U'�n��������mӌ��<�g�H���.�%�67�_><���r/� =�dً����[t޼1�sH�{09��r \��.�!CQ72�@�ǆ��H�]8��f�N k����sz�r�����dI3�[8|�xE}��������٫�w�����hA5Kg��hO���Tʬ�S�x�e�#`���m��gV�=0�|�H;x��]UشA�5��������p�sdn��-dN�	|`�C��'�/>0�(��F8��e���h?��SVQ]��m���8"��6���,$d���>��<d�`y������bsQ���	�8�@e%1��s1yk���3<�����4���M�v�?��V�t3�*5@؃F*KY��x�R5�:t�H���;^��q,�vw}�AV&A 4,j��S�A��j�*̇۩�η]�G�F3�`�x��ä���t���
8"���͟z�%�q�L�"��ؼ�RF�8W%�������A(��3dlF�b�~l�aj�E�ֽ�H<	�EuN�5$���H��<|eZ@��l2�K��O�<����iE/���¾�d[����������ҙg�o�Mͻ6=�ź�É�T���`
����~V2�4�,q�;��Z�L !���И��p��=���h�
�f��'�FY������£� �κo�5U��E����7�r��U/�O�WQ��=�����H��O�/�;�$_Oi��xl�5��o�)�mpDN��#���8,�Q}��bv�c[C��������P;02��]���D��b��~��Q	r������'��XR�_`B���e��g_B�Xox�.��Pe�X|��߿��;�8�ϸo��t�%�=cH�Z8u�����ƽ�8�}��>�a���{.+��n����<#�{?����ۄ��9E��,c�镅⎕�4{��� KfxC4�,���	��Zұp	�xI�����Xd���1f�>��C�H?�<e�s�a�{[n�]���F&��+ڹgPd M#�R�C���$��ղk�H�����&EtVE�+�@�l�N����:�E��q� �Ќ)�ļ���Umm!���4ew�0�K�X,�����y��Yȯoa���?\��O�y�m�(�'���A��Ģ\������?�&��N�PGW� -է��ڶ�Q�r��K���@ah:"�q2~\9�U�h��@��g'5m�5n�,ͳ�� M
]�Y��~Oܵ�K|a�J�C�5G6�IB��Is\��(h�ꨍM��.i敩�һQ�����b��F����Y*�0��Д�yN�����Ck�<~�C��]�y=:GA�#����v��cF�p��c���W!
�ؒ���X��C����z*� _�"��JVub/&��w�7*�L������ѯ���v��OˀY[[�����-���-ٙ���8@���__ �O�λ�y���qBe�ch%YҚ�&�\�5��˭��� d1�wr�,�R�|A�
F����:�7�Yn.3�	H�<k�d��Ӹ�~��2O��qf��{�&�d_�@��b���3'�����L)�DmCW�S;.����b���)�矯��?��4��	(�wz�Rq���	WMmo.���M~`��-���4$����̟|�����U1�9<��S�D�׸!�|� p� ?���g��X�.��K}|�[�
����k's�Gۅ�Ǌ��ո���%.�'��-$���vx�bJ�j��>�ר2�ŗF���l��Z�C��_-�:�+l�
�p_�5�_7^�*@DX�	%I|��:�P"��� �~ᑰD$q��(X�J�2̶����BuKV1/=A��YS�v�&9����ї��r�
|N3�|s9����w3)�����a�D����S0�5_K+Z�^�4� ~X�?Y�����@��#,Z��b��L��3yy��Ӆ�=�����ɐ������D\j�_��_��_�s��|��h  �:Ma�~���ܱah���q]�4%h^��P��l����A[S�� (�$��]{=�͇.�0ZE���{�Rd������٢�(� ��ɷet9�i�8�,���X�e��A$,��<�ڙ���xޘ�?�n�ם��t,Iq��|o���Z��7�zXv�;<,Yԯ�Ӭ�Ҵ��Ђm����������S=�J%��^���iM�.F�buVs��ղ�3f֧v�<=�K�T��t��~O0�F2vլG�0|�4=e�i�Xe�rkI���w򟖡��ӻ`� ��_��M�t4��ˍ��r��"���߹$�is&�n,ЂH��9�9<��C h���vib��,y�T�{�7m����1h���K�M�4L��8UNNVe�9R�u�݊�7�"Ϡ����xPu+�dJ'IG�5��-���{��46��?�d"*=UP�z�S� W� ��2�zO�kc��Ft�	`�*�����z����1�C+��7����ǆʖt�lt��UA3�/e��F�.#����uv�f@����f����c�E���U��� ���L}�c9W�?n������Ju@���d��~	{ &9��#���\~~'⬥�D|��e�����5�4�I�$(\���W/+f�R�"l��E_�׏J��^���3��X�E�4���i-����9'�����4 	��	v���[����/���0îp���x��ܐ�г6<�Z��/�x9��J�E�׽�<����~�4B�jye�A�+�`چ�7��Tg;`v!���߭0�p ��4;�7Ī��ѷmT��/�.y��d���'�l0r�1{��I ��͹�bP��RLT�l�`�Z���i�<Ԓ2�a��H�i���-�˄�:�M+���^F����{1<(����A�m��CZh8X�u��#�&�tQ|0��Is0�)|��oni��3��n���}>橈݋צ|�پ�kEz_�}�}���:%B���(�eڨ��[�>���|�-B�}�m'olX�!��;7$c�J�=\����c?�~�����>t�]�q�T�½w��DL����U��R��쮑�t��
����1,�r��B p��|i$&)}1 %����'ځ��EC'����#6]ͭ�W��u��V�6ҿ�V�4�����v;4�[�?-������$����sDN��v��W,����^���X,��9j�}�{�ı�{�ɚϔ@��?<%H���L�V�|��Pe��LQ���)���Ey�sG@K��y��A�R��T�0��)�r/�����g??X]��
�/^غ,���~��5��t��y���l�Ǌ��٨��#a�y�wЏ����(-�վ�o��pr�D�\z�%U[�	��0]�6K���{3t�_��KД]�� І>�Hjm�.�Zq���Ro:��~j-����oZaJ�K��� �a����I��*Q��y,�� i�R��&Å��ĜɄӼl�gO�JT/I��Q��W�����߻�.���65Y.����B��*� Eb;��_H7��4؟��ʔ��z��S�>��\���m�ݭ��Uྃ��Z@�&W�w��)�y�4ua>�m�����|B�Bk�� kz���&S��T]^��>���! mH���CNq+���������l�*}b�>53d�>��Z�y�<$�Dx~@�e�oR�J�����]	��[P�(�JZq�
[s�G�k��@k�`��!, T~�j�.��<{��ݟ��cf��0:��t�)D�
�������+2d�|BYx����܈^�� Z�A��p���)Ƕ�2[>��H���J�Y�^������n�dy7a��1�fz��O?t�2�P�㺓\9�\��8̐���Ko��ժ_���R[�H�$�ol/�t	�Y0tn����Һ�#�@��L�ؾt}p�D%���ʎ�����q b�p�X$p8"H�݌4�~�a�<�J���nZ��#r�Pd~��Ė�ױ$�77�!�k��e�P�b�V�9�����Kr�H�2�!��vͻAy�ܜeD��k�{*��j(�I_@����xe�F�`%��c��u�7c���>l�ӈ@*%}L�iT�5[��h��Қ�g{��wL Dk��q��l�}!��u����S�����Q-����`���ܰ#�\��s�.c�)����W��T|�C� ������1sl�������S��oѵK��M�<�q��8�ⱺ	���r�n�����Be����z�)0@�L����ڝ9���FE��.���̃��e�TQ�4�����żL�<�Q��zlW# �ZS1�d�i[��]?v�;�LR"s�.���&�\�(��H�疮ל�j� ���0���
�*��_��������H&��̰˥1�C' ����>���r��R32֒YG%0�[*�O�D�5�P���%�c{0���uC�h�;^!�iuL���16�ժ�Sz�ڬ�Xx!১d~���ַ��j'R��V���:�j(g�@}X]x��۶VG)m`���E��ƍ�m�T���
�=O�
��<�؇*�������d�(�n�P�r�䙮'kʂL+��c3:�q*V� �ߙ>X�w-�vwv5���i��7r�dS
c�EEj=>=��yH@�x5�l�������*8��}i鳅���1�"�,�3�N��$Ԍs��� ���312 w�q�KE���QKL�Р3.�#PVk����∏[3s�=�c%6�4C�fD !�F7 ������ss���$��5�Ƹj�����ޛ^s索�OPȹ�Y�淠4xQq�z�ٚM��\��%�`��"*e�>$�PR��YASţ� �Ň`���5�Q���(�Z���7bk�����$m�)�u���I:�f��A}T�ǒ��
,-�$A��*����A-���wX>9��r@R[e�Q���u�u��1��Loso�w׎>j8���%Gx8}xn�$��u˳�x�� �~R��.�������n�
J��W�#�R�K!d��Z��Z4Go -�Rά�bV3�{�޽  �䤤t����qcu�d�߬B "~�����Kb��ޢ�;���!U���ܶ��J%)�N�X�-�����x�Ktq����&|�~���uJ��9��,뤼B��f�j�I`�e0j8�KZ�9������8��p~I�+>Gt�[=�N�̺@�K����QE����̫t l�C2P={�x*:w��+B���a֎���&��)�y>X_:>_���a�F��v_�����uo-|00a[R���mk���w�[�(�8R���=U3bgǏ8d�	�!pDR"{f،�NJ�E,r���3n��*�A���� V���\ �uE��	V��Ξ��Zx��BO{|���a���)C�vE�����P!|�U��B��'T��xɕ�����ؿ�Rl���=��rI�)K?�B�n(*8�F�1A}y�Ѿ/��kҤ�:rjO� ���n�C�r��x֭A�������(ih�6<�����Y�<j0\=1�r�~�V47�_b��t�`�z�c�"=U�������h�g�)�L����6LN�r�r��
F(S��b	5l�.�O�fN���]�t�y�_;�q�q��f�жe'��Pa�����I^Hk+�|v[�j^E�����13��!Qt"�(��W9	h�k+ �s�qc���~G}����w�`�.>��1y��������%5�C��ry��Ĝ#��O
���R�����'�vW��6�����R�B�ә����F�å���{��e'5�jI�a�i)��7qQx(�˒�/�-cVm��P#UB�0}�G�S�@��y���*,Z q�ۧw�U2.����[C-"M�n����W7?���0�gI�p�qB����˄O��x�Z���t�~���.&���!��3<8�1m0����y9ɀ1�?�_y�W�q��B4i��@܉?�L��]Ν(֛�E�ߧ7o���-4}���Q�j�<ء��A�3珘��R�3��-����ȝW��p�ͨ٢��f�G+J���b}�'G��"�"C�C$���z�`U�]�� ��ab㸯z��|�}dM �>��x5��Y�!���<�6�7[}�mi&�+g��l B��
d�q����!A!��~$Qk��s~��@#Qj��Y��܃Z�8M�����5?��<��L]�br�*�s	�T�j0�M�A��������>cx���h���k�~u�o�k�}tQ��lg������,]Ѯܐ�����-�%y���.���GQ6hn����-ա�&J]��&1�E��8Y�gp�Gҳ	아ʞ(g�g_*�/{y�V��[2~j����E�[ ������,�}qͳuȕ�ij�]��ؽ
'jWv3�\HcVJ`�����|L�^�{��f��`~߇��G�ȃE�Q
T��2��Zƛ着����kw,�/���
����:F�.���+f����47¹R6��?�Q�~�%�[�r"��~9�3�w	.E���-���ޝ�S82ͧ	�!�ig�jCk� �� By�;�Z�M���;K������w2=n�|�?�х����0�#�z!�:���Ζ��⎁���`�mnn�2O�K��O"�QFe��tt�Ȼ��$���у��tx� 
��P\@����E*����*�z�n�����ǈ� ���*��TO"Mog6��T.W)�R��˯C��ĳ�N�V�ߑ=� �~�GⲄ_����<LW�	�X�(���v-�z����Cw�f�����h��/�\>$�h.n���Y�'����˺�Xҕ���n5fe$\D���|��a���>D�#���w�@���	��6�p	�w���j��y�Y �ŠR����ؓ���������H8�œ
H���:n����,VE=�Ov��<����K�~�H�
BI�$��}�j��'����ڹ�����<(��c.m��3��2J���ԨuY�85�Яl��&��qJ���\h��˞
Gy�8a׷b�'8]au���jzEN6�ޤ����f��q�k������w��ac;�b{�_��T�"���<��{��m�n-��r�E����\�����U풮�\�'$�Q����t��n��N#�Q(�PbL�S}џ@�6���A,#E&K��_�Zc��#�&�i���g(���M
˅x�8
`Mn4�G&�y���]�,���L�0��7G�tn�YM)�Kշ}Q�/��ø�H���E��ڨ�e�㚢�)`p�׊b)�5�;~�^�w|Uз-1~0/�SXVb���#(m\՜P�ti&y�f!��x�^�ev/���N�	�M�j �i�����i枖��p[9�B�t����:�{i���M�jz�v���T�l���2�~aÍ���,p�*BVb$6�Oޠ8��� � ������a�L12ۈ��f�e�p��ݠ�̓��
In���y�!�&b&/��d�F�8IC����F���M��F�^�J#�����u�Y��L*x���q�%5��n��"�E-(8���W��pe�sC�&�b~LK���p�F!�  Tm��rR�᎝Ƀ}�Խ�/�)j ��%B�M���аg�L2\m�`zwKn����2�ո�����L}B
���*�D��s@�-�9�TX	g��#LE���BA�ٸv-��o �'r��C�����Ԣn,A'�geb�� �G��֫��2��0�a��%7�Ki�{�(L_Sŀ�GB7FdL�F�MT�p���f+��b�g�����~��#$J�`�F�H��hYQMǹ��>���Ή�w|�s)f���?@�v��� ��`&��/U�5�`��F��弁?Q���A�|��evK�v�n��H�5�-��� �}�xiy���d���ڌ�"~#��0���s ����ߥ
Q�!J�4E�Z��ΖHFw/�vi=�_][��l�e,����n� ��y���Y���LR��Y��z��v:��ׅ�5��|=뫳\$WZ��@���
��v�+X<L:hX��n܂�}�nFX�r�b>�Eu�3E�@��[��N$���S���1�RCR �#ŜT��O-�5|�5�Ӯ�'OK"����*-m����1?@��4q_ ��Kֿe%ʐ�� |��U܊ǜ�8mT��)��!2��<Lm|2j�C�n�<��]ч��or�����<�x�[�N���ם���8�#�1ו���[J܂�|����Qo(�o6����	"���ѓF�+�ІM:��Ղ�(�T��.��B^F��r�&{	#��X���5��x4���+;���O�F�ԥ��tQ��~ mP೼�u���ɂs
�{�f���o�7�"��BQ���mi_h�����𜶏��%Iᮥ�����|�Cy|����?��x,NB���d��5�����z�.܁����r0����w#I� ����)�K��EE�kpis&�4���3�F9�:>�k�������Q�?�����p�J�N>|*�e��]�_$���������[1��g�Z��%���	/k}b�
�Z�����M��,j�4Y~K�g'�&V�4�9�m U$k�GA���<�wsz�?�6�{w���V�6������H߆
�d0L��Cɣ�]�6�~ݔ�]�)�{?��3��9�b`����0I+�����K9�O�lJ�՚!_c�=�s��Em��\�Z��-������dZ�*g �[����c��7+U:��t�ۛ\�4��*M���L�CU�q��<�:+5Y��F3w����]u�V0�_̀A&�5�16�VȬ�~��9��ڤ|S3�p�k�C��D.��WD�'��j�2�(߂�j"���=xe�V� ̕�l�SU��,�x8�Ȕ�6�����C�7/s)-�&Z���6�Uoĭ�K`��.bZ�7��������}���p�X���.'Xَ�x�ֈ�Yag�K��dh$!�h}�9�gà�!%�\NI�e��!p��g�4�v��Pu1��#����8;	��掦�AN5O�m�>��^��Q';��-�/*���6Q��q&��ܞ+��+J("�PJ�LO���Y���_���S�m]�8�/o�����}��3�x�{F�����KY�]��q�Vs7�fn$'��7�*���K⪏�tCE��F>E�U�"$��th��q�Ģ�����dUj.�ߢT�L>ntX����(���},���H�&�^aՎ��Χ�1㼉���R��{f�9��5�ku5<��$��|��]2_bD;���rQ�5
r��k��I�|c8,��?������ᶊ�o�CP�S�gw�+�ʱ�J^)�E��G�޸1�价ixI��"�q�9�rb�Q�d4&�"R仧>��W+K��8����> =�D 9�O�Z]R�l����O,c�E�vKw85��5
B����ν�.�'Q��~�妮+y�ԩZ� ���hN�\�����l}&z����"h�Sl/M����#6 '�e�{ހ�K RzJ�uo����	�_���b��X�����߾�]&	�~��D��jƷ?��FD�D-��&��.ۄ��-��O�
w��A ���^>.�e�qY;¤jL&��Rh,<~`]���	o�P��}f�<)�Ƽ7Z�ٛjA\s��.`V�����t~�p�-���Os?�0u{YY�=���|�N%WUG�.�p�+�*���}�Ȩ�)_��)|�.�����O��B��.�&�hRX����!������Q��'�io
�6�_֫�u��b�c9�c��=ح:4��;� �
�4w�O5��[��7��ῲS2P�&:`����Y�4X�dp���;d��&���Ӛ%�(�R0_|/-�6ɱ+8�n�;Hh�(%�M���Bb/F]�VY4��m�����Z�r{[���LR��kYNۯ/�Y.Y��kv"�����Ϝ�.>�YdMI2�;����
�0�|������y9d^s=���Xd���g5�}�t2�/b�^O���1�i����y�c[��RD9G�߭��c�B��[�j��좥��wk��A���77��\5� }������n-���[q�փ��٧�e��űv�D-��|��<��s�u4@�錰ZqX|5�����)?�cҝ��-[WE�����!7��!���d����N��m�`ط��OR�j:'�?�����ks��!�������?d���;0�h��@�.n(I�*��c��-$.�D���u�4�z�G�X@�y�u�a`�^�PV\���.�>'���Lx��p�͎>�2}����/����@�t���]>�|c��ٗ�bֶ]�t���d�I�b=ɍ.�B�Uc�|_�.(���h֟h��j�$_yJ�j�Ⱦ�-��X�۟8��y�{=Ɏq�J�/לMl��
�����l��[����A�E���5YV��L��(��G��z�FA���� �,�O��/%�'�&Ùg�^�7m����@�L���*���8^�Z�l�A����/�U:q�ۈ��^�����|�KL2T���7$���]���6_ �8��ӊ1¼���	 �?�@���ǔ�f�[ez���	�����e~zb�-�Q�X)�3MuZ���n��ihk.=�W,�� ��ҫ�R܄=����cdĺ�զ�,�aj;�d�#阊Ckw����0��U죾ω�=��Y���9���|��mK��HȢ�m�����|pGf��7'���%B_/���j��@�����#�R�>U�p ��h�ϐ_�n%�ئ�>�֚�����fTݔ,�����jm|7'�\�Y��ɥ��%[�� I��#��O@�I`���;?�]%�6���A�ֲy��4��?��G�g���Yg.ט�K-�L��v¹��F}<����z?�]��LAzk+*~��Ju�B� �<�8���Q�}����m�:Uq���L0;J�ݩ4����5����鬐e�{u�QԔA�3Ô'�VT�Q�����>��Ԩ�⚁|�E�S�7�\;r��n�{
0�		hTy"���c,# �����b	��'�SE�_�GO`ZvH.}�t	�}�75�,���4�HD?Ǔ�Rң��[�~���>k3 sC�F㇙KR��'^�ŀ��dp���>��P����p3=A���dg�Ec�� 8r����c��?�\�]���a{c?}�z^w�"Db�u��yøi	�-����k�װ>M�ٵo�I8a���[�0d����˞�n-��d�x�|03QZ)����m #���������<:]6��Fs��'N�Xھ<�mQ�0뛌������"����|�
��w�p�r埭"�7�_o�+$׹�oMm��M^�{Ia���⊎����P��W�]]�dV��+ &�w�6Ɵ�0Mi��N1d��,��̷���`�nczH
�On����l>z)�*X�u�/� qU%M|�u��p�@/�((:k9��Sm���֐�#�m���4�K�*'s�����`j����/���@���ք[��-����S���b,�!���^7�+I�F�"87?�[�d�
�Q�i�y&6�������i�%��I�ry_W�����=�Z+Vا���!�Zd��5;W�W]q*����~:i�ņK�;5�j�o˽�wKn� �gX�݉?�Z4��_�Y��N�	E^D��i����r���������g1�H$�ڌ�+����"}+� �_�JK���7�u� R�a��e����R�4�4�WD��s9�b�O"珬aoA�puA��}V���Qu��e�������+vbz��>0T*��3�1_g2�f(�*ĔX��RM~>^f�:��A1Xp�3v_��#_o�q	����l%�����tVgS��v�ǝ��ad,�g]�r*K	t�����a��O@y��`�yb�P����s���E��R#lR�8��Q(/�t�Wq��o�l��pߟ�,w=�[�Q0���y~�WN��F0�״]^ru�S9��-$�9A9ֶ�t關=������Α��!���������Y���=�;���ܚ��`�'7��]y����K�R�6S�d�hw�L������GH���dt-���~t�������<ٔ���ן�&ߡ��͔����_p�~MY�E hn���y�P���lK�����r$�c^���B�	B�e��C����;��B�g��N��"XeB��������3���,,tK�!��Z��,ԅT�A�h�R�M��4~\{�kj�1;4b0�J�C�孷t��'��pȦ
Q:�j̓�!�/]>�r]�A��SG�q�L!�W�N�ʠ�� �d�"�Čب�_��L�>����3��:��ЌP�?��P:�=��x�H�������G�_�Et����9u���eE���9�aӊt��2Hd�#ɷ�I)D����Ӥ�S������'j�rcu����*�%X��p4$]:H��)�:��>n�O��,r�v!v�c��Z�HQPw8a��>y�_�˵^�I8/�� Qgu}�5]��x�9���Y�^he�k�\�ޯ=�5��
z#�ltu�/*wG�.D#g~�x�"����oS�\�"�A٨1�K<n�e;�`��D���J�ٟ&-䎩kn���a��L&�(i��)�D Yw���`dfζ3��g���:�����q��4j*�����ds�i�e���:'@4C��6��y��N�ED�D���YX�ī�JR3��4����*(�JԤp�Z2��9��5��-ڂ`2��^��a2LN؛C!�J�� �RH�G�:ɀ�ݾTn3;��lQ
�8?N�bf�6{o�;��Wɼ�_�dO<���#ջ�3��WpUd��@T�OR*z���S\f���e�8	��0,�)s�m,��q'��^<��=8���R�����$�(��_?%�� :綟h����D2�F{]��߽g�g�;���-�4�-�L�~6o�J�Ŗ~CZj�K{x��=P���Efȱ@������;1i�3>�쬜�H����b(Щ7X,>�%ܶ<�C��ޢ*���ceC[:���BxA���&R�xo�L��f�N���`�5��%FY�-}��q�zs:��Q����Dq�,鎼1%��3�V6"��L�Rt:v�g��m� &�)�����Pk\����䱒Յ��&�n���瀄��~5���V
ݛ|�ag�ʗ��K��5�}�(���ϕ�����F����8p��t��f�J��Ъ�.d$?A:��~N����tnr�6��(��g^���^�!s���� �a�²,��u�i*M����v��0��`wu>W.h�J}�--�GDb��6B�YbJ^ծn)��O�Z'�r"zr�RS��^���bzy+�����������f��[�Zǅ���7����O�H}��<8�υ�����z h�I�oX������Xx+�ѥ���
id5_6Pc�Rl;��\�ߎr	ی��.%E��:���{�kF��Vtc(�EҠ��|�_׎h�Zl�cN���/9>���|4ǖ�ƺS��#2ı���7Pt������J�S%�,M[���@�*!w�g��΄�%.aҴ?fT�J�P�]}�n�`�������ᛤS.����Q43�-�g/�~2����3��+��^�Љ�J}2w�/.2%�y��/�Y�O�gk�;`Y��rS����&X4���ln�Z2:�d��le�7������,4��k@ȩ��^����!Y�����i�F��-���j�5}	���B����6�k��e
���߻��c������C"��3@���Ľ.̀%5���zͣ�+A��TQE�E��H���N��|�L]ź A��ە�kZ��IΟ1�1s.y І��GQ���]�LQ����#`J0.�m�)׏Ja\@�D*���?R���c�25DǑ{4��y���='Y؁5��g���M�K���3�qh�;�1��
�W���!��Zg��n���'�����爜�+ -(q��f�P����_^��im�p�5A��UA�$+�B����ҊwLl�vjG��L1h�1�|N�}��̂�@��k��-/��L��`��^g̤
�O�-%n��r��bѷs,V�l��/`�Hi-@N^�j	�x��Bb�nZ��6�vl�i$(�n�C�1�_+D�����!Y�?��.\Z��]@B�,�$-s�x7E�U���p��L&N�� /N��e/�Ub�1/=VM�iaD���짆=ϊ�f�Xc��}ɝ�U�o���l�;�ܦ�S2*c*�k �gd�f����/yK��M�r���WmgM2�	P)��Yz`&"$n+��8�%��W5��@c�%��d,�L�E�.�D \ �+���}�� 
|A-����5�c׭)����)^u���G2�f��.u��n�ʚ�&ܶ8����$�N;��;o����5s��^�s�`�.Q�gX`����kя�
��x��xCمuH��^��)
��D=?z�x���"��UitoT)7�DO �'�OՆ�<��(>�8V�����e-$Ue�=G��O�J�hP	%B�tȍNTvL���t@e�E��ز4(���c.�t��ӏ��/Y^Ci��>N��S�R2:���� �|�y]�O��w��gCM�D^?����A��D��i� >ŵ��0�x@f_@zJh8�:����p��D!3�-�H�w�:s��>h���,�g�S=1`�?Tt��:.�|dt,}�.j�SP�3�]���g���N�V��䞇G����z?*f��,^�� ���3�527�G�QWf���p�C0���^O�R3�=̐�#/lԡC���Ļ� �S��<.!QmL��[ރ$����ȼg���i��U��T�Tu�t[�n#�vG`��H�k\���)C�����A�E�٨��x3}�e�NY��}^�}��D�0�I���"�*;6��;f�����"=��7a�e��L�x/��kU�P}ƽ�5�äO�n�*�uO_�p�"�T&�~��>���u^i�	1�l[����>Cj�(����N$E���&q�I��Ζ^�5.����"�붷ecB���u�� ��u����ŧ
���F$ДR�\ؔz-%"��ѫ���5c��h�,�Ӳy�t�&�e
�ٷ֠�o����"\z�֊�q�s���1��.��u��X���f�)���E۾5>P�sϮ�
_��C୴{N�&[�����!����� �g�f�O�n���,��)z6��3@j1�6�S�]�R��K���0�?�2H�o�ղ ;�^�l�*@W�r��A�G��ǫ��_Rj)�NH�u��9�\��q�S�]C���M���of��_����3��{!)V�-
���e�2��̎�:7L�[,�r��#Zٸ<�M�XRv˝;i�#�N�L��ۚu���A���W����eμ�+>|���$9� %:�&���qt�E�U�C-�?T���.{� �����k'�z�s�63>@t�7���3(i��B����j�I��������I;�Nȉp튧=��U�b	ˡ�3�p���-����-�� �q���g>	
{5ލx �$4/�_�x�(L�>﹡0U�A���S��a�	�pͭ�`���0|��� ��^
:�������A1N]){�|Cm�i֣9|�M�-�	����MZ��ļ��7Bfz|�Dg&ZF��ׇw�����5]s�T���/L ��+?�wx��ST��7�7�pc�<�W�2i���ώ�'�ܰt��P�yR�����r�Ğ?UUQ�ⷪ����8�^o=�������q�����'`yבּ�mU�����K]�uy���K!ؚϾ�&���ǯppZb󊕊�ķ�?�;��7���_���}�JDN 2�oȵː�Z&4����E������{�kGH��s�d(sl�#��i�q������r�_�?a�v�5A��.TҌ���<]�,�_I��ʪt]�I���, ������H0$)�D��"�A��&D��NM��)b���w �Z9������
�3�7��@r�*�7%cM� �U\�eX�RFc�?l=�>�ǻ).΢g��N¬ �=OV����"^��w�9�G�K3i�w]������B��MTC�ݖ��.�}>�m����*�N�M���R�-�CW�y��ˋ�,��4W�@W���$�h�����w��*g��*~���ﶸa��S;��r692�d%����L��U~P��R��e]����!뾼�83� �|��8�k��dL��l?A-�k�a��[��c�����t�|�>�#���!�S>�+K;D�
�WP{vUx� ��o[ի���YG(!-R����g�lG��*��	��a&>xM	�=š;
��V���-^���Y�Tj�#!*y�\<St���s��i��i�6��0X+i���4&��=�H��ۑ��@ ~��.Hto~���FA尒w2>�P���rV"w�N��(��6��y_/H��w���X�L
�N#0&nNx&˒3E�`@b�����EHvd��0D?,�۾2�'Q
�C`�"SQ�XI7Ƶ��4���}k�^��:�;\-��?�@��=(}�-���/[��4يQd�69�㖴԰��/�^���Ӂ�
�_KEH_J�ʞ�V=d�9GBK����?��0�KZnбɷq�;�(�hå���mOq�PP#��M!��?����sH
#���,V`D����2�zo�X�v�v�/�N�i���p������ν�R�&&1�N�c�˖5z9d�YK�E�e���fnow��{Q��|4�ˋ��/�^	w�ڜm�I6�j��ϦC��-E���ߙ��_Fɷ�>�]�ۺ��;�fD$���M��y����:�%���J��{�T�A��t���1k �Nfx�NO�+=���C�C���%@H婋�
M�u�Np�j>"��٭<Cfb��!��4s�ȧ��؜�������I�E�J4�e&�F��������@t|j�א��~�~t���̯��Z���
�,�&<�=4�B�����6 H"C�d���	��]��􈦔t�f�#�C�cy]TVOT��2�P��yr)g�5)���i׉����枹�S�q�YWE�]F�x���]�r	W�8�f�����z�eh�7�^�k���<pdF'o��������ۅ<T��{P�!�-�O[���"-a�u�4/aLȾ a4&��x��e?�B���y��.�E�Y��9릃����C<�~W��}ֻ���-&F+�r��&K�^S�A��}���r�{J� k*��65�tt��h���G0O�xҖ���Z���ʑ��u�����\�>g���zC؏���
�~(��^���-�#>���K1��3�>x
7)�3�'���*���V{�.Y�CQ=�(���$�c����.�[�c"��-P�m��;�)��R�X���t�D+�~�p� B}I�� ��φ��G��@}�-�`��-�G��k�:��Frx��D�����"��@s�6D�~�d�4��VʉPu/�y�"+MZ+U�{�?O%�)B� u��v�{x�S�����-/ۥ�>�2���#��WDt�I��e�C�EY�\���g�c> I��}��)�hG���7��v��@�w��ޡVbx�n�џ��s�1!��~oq�-mgo��
hH e>b�֭���h�:ߛ��1xo�1�!�Bdvݦ���C�T�������@#&qC�l�Y�j�;Ss�ډե��H��e��yD�{	��-��<Z+y�40���N������^�i���f��_�juM����APf ��ʳXfn�=�Ж㢌�fh����=�k�_ ]��?ј���|Μ�7=�`q�3]+����xi����6��E	��.t8/���P��{�7Iй�iN�[o��c��Z�TE�4MB/�����#���\�&��8����t��cګ���%!�Z�������	) ���W�D$��<za8ʒ��'�{#�Uz2kB�/%���������x��w�<�㍏��9�,e+Ϣ��|�&�z%�1�u�v��� �'^a�e٫�7���o�@��=�oU��KF6��7�~wb���Ő���R|�6��Ŀ��Uw����_�@�=��p���i��A
]��d�I(����0�9�V=>��|z���N��S��"R#���w`�1*��"��H���º�� DBH�:��@x' v��nc:���N�G����!v�٤�pbF	=�?T�2j��O�����A�&G+]��#�`��~�K8�g�����4��f(�j�@RAϏ�����YHc^�J7ֈȉ�Z�9ޮe�k�+99�Z�T�{̅��H��(����퐒7"B%����V��Ī�+�e�kџB��ܔu���VՓ��	I�~�B߆���
���j���g�(@���>y�B)ß�q_I��[�KWuŀ����R��g�cb�P����Y@M8f�|P�)X�@�� >d� Tȟ��w�4j�Qq� ����P������`����}�[��nn���m�/$:���&s��K�j��P(Ϭ�Z��0j��C��a��2�p����H��H��l��v��1OA�,�z��g��*�B/��<�EQ�^���kC�
����O���w��!h��iz̔ء����J�o�_�J�����X4p�����|Y�E�9����2��֤ײ݃I=^�����1Ž��y�d����p$-���P�d�m�{?D�&o����<�����w��/!��GH5ű��?�2�9f�DO��h��U2�v�����B��m�D�A�vjQR[z�,O!�B3vȨCYZ�z��kÑ�LO�F�ܽ�L4��m��.��J��'�V�����#[䂫,�����a"T;r`��=Jr�}'��N t�=�� G�>|@�j�u�3 �C��C"�%��z�P������M�"N��Kg��\)���*�_U�^�;Z�}�e����W�Ue�Ͼ7�n�$ȷwE�T�98��N_�̿\��ndlT��!��C�y�J��,Z��zUkn
��9=ǫ��~Μ_a�u�i�U�t+8��#��~&X�k3Ex1a�i�s���!i>��&��r=��m��J��yβ���RQTu�6�탏�O����8����~�$ ��Ap��jι�}üH,d�ޱ���IV���+1e��X�����^7>����O���_�D��}��[P�ǅK���@4Q�v-��4 B�a�udz(�ᔜc��#DZ��0�7�[R4u6v�������H_�:Xu)�d)Q�5VEφ�.ӣ����G_`��M`_+�#��JK��S.1��B� �[=�+���0ǬԽF h4�ؾ�wh����ԗX�\e����tB���/��y<����Q����k4���}T��@G����S�hp?�����Tp�����͚�����j/X<�Ro�n�
[�-��kF���&d������M�0��=��y
�z����:ꪖ�8��\R��+�v�1�)O�D���`=�D�O��U���5�C��a�ǡ�ګL�%�n\�ԍ;������,�W4`vC{�>;��x��X��R���'����OqƘ1�S-\9�o#�f���I����(S��D\����@��}���-u}ۣ�z�+葫i���`�#��;h�3ϛ�L^�TN���������
P�)��Ʀ��t&Uei��	NR+��̍�g��O��A$�a$tȡ�U��ޔ���=9����*M���BGnx�I;�T,����Ԋjgђ�m$�:~.��#��� ���v�tۥ��׶���Jd�4d�,��t;"���.��^I>�Bi�3)��1T��s=�*�^��?RF�F9�GA�Q�h�0YV�۲T���(8�`m�4���ʪ���i|m�=B��Y�����JVS-�.���1�4�?���9�N��Fu=��Ҋ ��2��2OI3Ź@�S}�����G��f]����
�
���6>���g����RHXz6�gGk�6��X��%X�[V˔T񷑠0hP��h�4lͽ�k"��b��ru��Yw5@��2�b���g�����[����zz���v��?��:��4K�WY[���u����,�;�L�"d����,��Ӳ�B���j_�f�D]Oy� �l��dF�;��	/���Hvc�4�������J[��B9v�Dyk�����!*1b�%A���W"5�����	�hmEZt������4�3�q�"%���64�6@���&�W�M�Q��a���B�ah�"�'8�w�PX��C����NHq��j��) ��q���(NfLj�sK-_�C�8Y/�]��
�M�J��ӠoQ(��
SM��{H?r����ݬ��S��Lu���K�?�d0Fo_�n��
�H���ۍ�1BӬ�v��4�D�Z���aYt~U�ލ�ѯl�Qs���sz��5��������Q�.�&`�KQؖz���'������,Qy�_�0#־�^�qҘ�b^���é�X��<S[�W�5�@�����R�zc�S�K g���������$�3��T��B �BesC�aAȿ妉��Mrc�2�H�*U�k�?y��l�zۡy��8w�f�L������:���[��5���t�Z��e{ghuoJ���6@\u��/�>/@�j�R+��,`v,�W_Q�
_��V}�-��7�Z�ɇ��Y�͂M������I���X�Q����:�v"���F+vF�a�}��;n��Zs9D[?�KQD���i06��i�'}խ���'�:GY���E��!��#��r�N�����h!P��T���ۆhX���J*�9|qRX�=x�,#����g+����ihb�����bR
P��d�M(�e�9_�������G	�J��(�jtTH��"��8*m/�dO�����m7f}$��\�$�Is���g|΢h&]��D�L,R���Nz��|�p�T-�i�	S��i�@oh�)g��-��F��`�Q�e�i��^還�w���"�u?f���ds?�uC��VaHUy�{���tW��$�j�#׽���t]x=���|��Ty���h��S���yW"0���ܯF^�zDo�����x������%Q���J1�j[����\�DF�g$�m&�g*�4hy4�db�ԗ���-���%P}$ģR�	��B2K���>��*�߶p�7��6R5X/�6�ӿL_�mg'�AA勶�M�G{�����w�oԲ.=~�MF�jG�۴t nO�뚰��K2�}�B0��q��:� /<)B�[�S3#!%��A��g������_L�ծo?ue}nO�B}��x��nM*0k�az.\�G�'_ ��&�lǾ����	��ыF� GE�e������h��K��i9ڝZ�uVu��e���Hv������Lg�x:��>Xb#�%���-il%�� �ʭB�KK���*��6�? &�^�!P�*?QP ���V_^_Г_�n�ԥ�h��<2�Q�s��=�$��zAnal���� �S���y�:Wz�dO���>�S^��A�2�B$b�<P�˹\�HTD��|���a�}R��1|�!���=.!<3�7hE�� �R�"��ľ��S��V�iK��*�Xl��� tl�v�Iù�ˏ���Lȕ�������9U��<c8v�����usy���W:։�� �ap�*$�/�ѐ�{��kz��`��>}q�Ï���\qx�m5�\�7���b�sZŨ��;�r25�ZK����6Ṧ�/@膘vI������nJ�II�1k�N͉_��D*�L�����$CB���Hz��`�;�z}��0J��� �R�*|$f��S��؉�R�A>�5S��k�Q<` ���U&܏}	�lm֭�ȡ%#��"��Jʕ4��4��_�B�$�����rOA
����1a0����[K���b`�M��n��U�����i��� z�%��i�*��:�L~�i�O�E���G*d
u<I�Ds���S�IO!<pK�{�����o�,�V�+Y)��.��S*�]ΩH2U���h���s��EkN09�)Ucn��-֞n��Wp�F�eg����D�S��������}��X�.YR7�Ծ�����~� |Y�#c�����҈]�O=�[X�h�Q>w��?���M��hY��P���y��G5Xc�t���M:pZ���~��C�.-��Sj��~`���G0�5�E9��4�c�ө�a&L��]&��_Ղ��V�~�'�s~A��H�י�?�0��+RXz�(�"9����;��i2����Y|�m���+Z��j7���5Ph^ΘW?J2��(�/ɜw7�v��9_����9�R:�λg�V"]skD��Ը��pQ���)�n��1OE�0��/���d�*S��]�(1Kӧ�WT��5EW����v ���'E�;iPI�B-��v�����^�v�伧�4n���B��� �+e��I΍���S�V��mj����*8����K
ĳ7��;HpZ��b���145K�B��p0�t�%uɑ�n�����#����Z`��Hs�� �|!�������*4s�j�ϝ{��dI6&ǰ��O��ު��fݘ���6�2���53�F&���Q��s���5��	���y���}c����4�:! |ym���%�1��5
���jVa^�}����a��f�����puP�mկ���.w�`y�6G	}9lª2(s�d�\���T�H�ҁ7��&{�y9���H���I]Q����l%ee��
��?��H���p1|"vUsʴ��fk9_KF$�^��S�z�W�J�)M���7HW��K�he��ze����e��7`GM� ӑ%����2hH��q_��rb0p.�#4�Nf-USAY�c(�k��)S����A��Yy.	�R��.-{=� Um�m�����'�A�L3�As�!g��wq��Ǽ+�R��Z�N�[d�k�{e,�w��w��L��� ���jF_Y�"�DL��7��yJ�o���N"|ْ��uĂ�⍎��ҷ*j���{JY�_�+'��wrփ˛*Ao�io
�#\4�.��Nh}�(�G�S�����~�",�^7�g ޤ���1�X���B�|(S�F���Ǡ,�k;zp,F���uD�d��������"l�mF�3���C��r�"q^��� �������ܙ�Nv-؍��"��(4�j��C�~g�}��ĩ@�Ǭ)�%�)ld`�i[8�C���)��|��!�_n�YPdN�K��G}'��e�L8kO�s���ACF���3y�2�L���_�JA"+�(�Q_o�=�#�[iho�}ڸ�G���rο&���/���"z�RUU��й�Gg���>&l���o͡ԷD�a�H޾�b���;���e�G�t,ʄ���?��a����n�48�(�v��L&Z|�6�b^��(zr��k��Ke/�B{�` �Rm�ēHu
NsN��g$�_nc�%j=�Ed<rR�)H���A�89��`3�I.~� I���������S"�cR܏KK��,��)�C��������Գ���KH������u��FX-�VU"U��$����;��Djt��������8E�����2���n_��Q�[PQ3,Ng9�{�&F�wiW� f0H] ���!�a�o\���^c٬����(�`&k�X�\2;$�rR�1.�p��|��'�8Ս�U|-)���5"� ���
+��@�bk�,Wŀ�~x�����G����l팥�I&)h�E��^H��r����LENفRM�������\��3B>��2l��1t �wK���s�S��0��T2,��;Z9�Wn>1
���w�a-:Dpi�+֫&�S=7���:��]�Ŷ��$��&�I��g��3�=6�Q&g}�n;"����^UU��u<�a�-&��Rt m��Fm�Ƨ~S�6}�KQ�r�����;�hT��G��qLs��#F�l�'��d)��tS5(�L�c�l�TD�D�sF
h9�,�7�,�N��rFA�|�]��.��'�E:8�?�7�V4>�v��P9���x[��MZ�N�F�J�����-Jx!	H�lBz5<��KQy2��Ht��N֔s (�s���Y�sn�1>3D
i
](��nXV�g��0�4}���ʊ�����-�:�g�'�-�N�v�-�����I,Y=��A���@���n�%�i�Fk��g��(d�τ��>ڌv%+�����N�PpNiV|ڷ��։6]����mW�K�7�"4y6(W�$���R��mue�R����S���ʻ��d��q�Ȃ��
�@;�
�KGs�=@�SZb��.��W��ԅ�+T�������n^�m��a@�4�M��  _����td@���u�*a�/�KW�x�LS��a^zj�j;_�����skx�d��2��������b�Ee�XB���. y�
8T�W��)��s4�ٚT�͈�/�O���6��:��o�r�?T�p� ���g�Q�͟�>�'O���N���+u����ӥ�/�w�'i�2/��r��ם�&0���}���Ǐ����b��y)���79S�d8�d�w� �N��8����و�V_�G��)7�O�<ݍ;�&U}ߦ~���5��7,�c����������� �w��z�r��x��U7�0�����D�R����E$ʽ5u�����S�z�P�F����F� 77Jɚ��]607�1m�x`C��b�5}ú�Rm�TX�AL��B��s�1H�S��KUK�߆}E��5%���`=�",hF�SV�2S��C2�;��뼉Ƅ����-��G�'^Q_(a�[}�������|8����dc��	��fDV>H6�{|�� r���S��C]�5;�d���6R��
�����j��ɓMY�p-o�
A1�u�	�s_g�-�$V��1eκ������ ����s�P��<MY���oM�ח���6P�1�a%?��B�rC���ۼ��A�E��Ԛu ]&CVǬ銠Nn�l�t#b�V$K�4l��]ITё�q�����w�VIY�U�"�NI�D����gX�A��M69��"~�o!Y$���,Ls�H�����QG��Za��9|^ѐ�*LE����S��tG ��ejnj�1���q)cXn�Z�,���]`j"7�����(�Fo����,�Sl�Q����f��]ap����}\��K�O���x�觯�,�8���%�/8�e:K) \3@����� �D�c5N\Qm�e舼I�s��Mgf��b��(>	�[�9�w�UIugj9p�(g�5���#j��X�W�/�'���gB�;e���>�����;ɡ���S���{a� {�va��$��"n� x�}+����M�r~�e~X,3�}����IJ�쥹���*B����y���]�Z�h&;�'|_H��4��N�?�@:L<B��}�_�hE.u�c�*tB���q ���)KC`�.��16/�9,'�O=%n�&�x+��!m��CDY1GD��{h�i�L��Ix�8�q:,��$��m������h ���H���UƑ���S���r��'.� �~�ی�n��Y3\-gg�k�J<`吳��bk��M�~J}��%�����X���|**7;f�V�¹�JP���mﺘP=�L���hu~�B�9ӻ2�c���(�Q��p��M������ �|��-�-M�H�^����i��+Pz��2�
-������i��!�!"c(/�b�iP܎�M� >��J��0����8�]�[@_�Ȯ��(-!�`�2��g�	�
��e���ovKi��Z��y,2�$����)��@��h���R�����p�X�Hu	�A7|�����+���k����=�-Tp'���?7v[�z׆l?V�8'O���ʑCd�Ruc�etFT�0���+���R����tRc�O��@�qs�w4�^�Wk�������8�S{� ���I������
�/��B2��ڙ"�lU��uM�k��M�}Y�����G��T�Y�Տ0�U�H���ڴ�d��b-� ����3�\70a$Mϳ���Q\��sO����s�0�:s���-yx��vk�ȉ�cQ�~;�ڨ�:�u`C8[����]*+�9c��J������~cS��~�̼���o sWSD�	/��X���e��l+�Dl���@���K��q���<'F ��2M�ʰ�����mܶ�ܾ��Jj�k���';Tw>�g�T��u�||��ٕ�M�a��[��@a,���l������%�̳,"��2S�����9
c)Ђ���"��xI��	���=ejH�ƃԐ��}U*�'101����U��.�9�'���t�!\_��4Ly�[!B�SS��A�L�_0 ��17�*(a�q��w���*DMO8��'aϫ챉=w͏<�gf�G�	�4*
�]s�J�h����f?A��1��,�QHI�L�ąi-p[��n)����yU_��M���s5�ٳ��Ƽe��s�pE�s�gH?L�Mb_���Zg�����M�a���)OG��L3P�c��̱��e9zvS+7�R*4\�,u��#�Ν
�^$
���{��z�N/2p�?��L8����>�{.׎��4�W/��|<#r]���g�������_ڨ�m��hU�4{d:c` ��f��U�Y�՟���֌zu�A������2D�ɓ�RS������:��}�@���t�}��xp:�� ��=���7����QZi��g5ú��(�H_{ly������ hğz��_,@��W����SY:���'����S����N[yi$D�ﴏ$��ϭ(�#;�[�F�W�p�����7(~��t�S�0J7�B��<[ܝ^X�	�M>������,o�`gQjB{DC���јG\?���P���$���j6+Lղ+���E
e�.��1� �d���]Z�,�c;�9��g�>�~;�L����L_���AKeug���*�H��[�DlE8d���aq����\�GK��ma��e��¢ô5h�2R򉟜��`�ɂ#'(�����4,��p+����$@�
�<�,{�^ �à�4k.Q��=dU�]^��5���,V�N �䮓m����8�u>�����[1��&�X���zI�W��9-�@r�TdԚpR�EC�抵��E0��B'���Po��:?VK���0�6��*lM/�G�ml`��bI�N�>��5Va���A:�K�p=�f'�1�[q�H���K��D���z�P�2�8o 
"�roT�Rx���m���ֿp�w�s�\n�%��ֽJ7�98�$
��s�+.��bF�����Q�A+�v�z`�݌I�N��W��P���/Z6��3���rz3=�5�#����r�"�����״���L��loC�9��KP�Q��n?�\�곭�o袓=���=x�����>���П��w�X��� 8Ky�8a����j�Q0z���7����}$��$������{īA������,��p��t*�xh+�Y��}�������Q�"Z4o�����1I$�|eU>zP�a�CZg�a�����2	�Y]�.�c�'O��L�[~���'^1
E)0�9��KCu*opmmL��g���3<�-�������5�L����O��P�{��iPl�?�;Q��,�@���Pzaec���p<5x?�'Y��<���w
��]Э�[e�J�b�Ɓ����;��Ê��#w��կ��0Hw1�f<D/��l��q�~���@$f(6���V�˵�sY�o��tPv�_/����w�0�g
��QH�i
$�����@͔>/����h�iP�:�'!��� �Iύ!ҙ�_�Gw(na{��%y_S5ص�c���U�������[m�a�yKH�s�L���		���$�8GT=(��*�r?z�u�7UQ�-$_6��7�0��ޅ���1�*�"_N.�dzϳV ��2���Va�~D�O��3�te��r�U�12P���-5�G�)����C�(�?�1�Bx��M�^�;d���*+q�\�m2��4��b��Aټ�Yw���+
�2F!*4�Ȯ5zXUzf���m�: ����O�jo����&C���4��1�B-~]�=�,X�@?�+�W�	R���ڽ���c���?���x6@*H���
#��h$�Bd���D���O���qé ���-�B��)���',�C}�~:�Ĺ���6�R�w.�!�b�L�p�2��v	xfط��īR$��� u���,;����tv�U[A�r8��`�c��2jG���(\�o�SŔ
-K��V@�K9�5ERP�߶ ���`�9���O���a@�����)v ��f�g�b����j�p��Va�`(��D�j�>*2�#��%O���;p��c�P�""�\r�@F�ƽ�,H<O7>��G����%��C���}�K��j&��W�Y��11-��H�x���l�A1�5�@�H��D��*d%����9��!�� ���¦�d+�kP\������8�5e 
����:Yl]dg�W؃4.{(Lۼ}܌N��a�]&SF�q _~��D�z��ý�=y�<{��=�@�:9�0J��Oh�$�oOKuT���K��Շ#�K*R���+�ѡ��Peq�H�~s-3��d��/��t�0���I�q
W�H��{����R�v�4���r��ؖx/TE[��[!�#QM��S�B�]�a�/�˥��L�1�j��� c����Ue;�5����p�����8��"`�!�˗�T�Ŧ��s�;�/�>��%�a�
��T/l�.���v�]�<Z�Y_kF���<�Gk�%<�	Mm��?�K��"
�hO��p߼�7S.1?�z���@t���Էw}V(¥�*#	s'(V$�o8�.&�0e��h���u�|�/�Bs��fwY���.��˧]�]�t�l&�B��Rrw�l�g'�H�h`�5���Ň���t
��S�_ɜB���q%�b��ޕ�ѐSI�UWZ�\ �MK�
M�~.K��q�cѵ{��¢��ȓ�b�e$�y��2HF''���G�����0hK�J-���+�%��|�?X#�kT�oɹ㜢�.W�\��AK���YU��y��jov�-�����5��C�P!��Y��a�nO�h-#η`_�Ns�Ę6���9��W"J+�T���+�=��V.`�C8ߚߪ�!�����|�t,X�T�ڏ����L��d�����ze��b5�|����?Qay�n�J���ZT����wĿ�׈q�?�Y*�R�ddX ����J��Q�[<B��a�i���8=�S�?��k���.�B�����0ֻt��B�3�z��0Ϣ��sqJ����A�	̨۟aq]�;��XG$�.�Ж���1�],W����4�j�7��ϓ�mT;�$��P�`��,���P�Jq��l����l�� P��M��P�;`�+!7{1���=�����t������%��R���]�𭪘�l4<\$o��o��1�3@o�)W#��	���t+~���P�I/�4R,����vj�-7���|%:E�3�y�m�*G���\�c{N(����Zw%!��Q^���"�ӎېlڋ��R��]�EZ��3~��T�[pR���H��VAĒ��Wl���S�k�� �Q����'w�s���_���ۧ�~�����a�1@��'�,(>�yQ��6��h��l�o�uu	�)�n)��<7g��d�m$PFF��{�j�S&�����nI��\�,�Y���*���U�G_z�s���?�ӝ������2zh��@��B��*�4��}Cp�������a�S��=>1�H�L9���\��}/��kV��kn�`�G#�~ QT8^�|����@��*R��"%�%�&�9w�J�����bE��^���[0ό
��g�b$�j���ݨ�Lk"�{n��0�HlT����t����qBo��t�ұ��u��y��S+�@��i�)�۬"ڹƋ��݀N�3��ǀ��]��|z ��,�Mq�	TJ#�DBn<�>*�ߴ�&����O�L�I_�5�!��s5IPEb-�����c(�R�_Vbv��ޒ����m��s�x�Q���S������Q�4�m]b*�aŴz�-�U�K��<b�F��ʟ�����H߂�O��R	�=[Щ ����)�������Ң{�u;���d�m=[�Z����X���3�[r�1^�j��A�o���?"
���z��K8F��U�L9������\4Jx3���]�'�����&�/�Ƚ4�<W
Q�ך�^'�9k�)Ϧ<�p��T}���ӈ$�1�,G��s�����󛘶��s�Ν�a�{e���?�ﶣˣ��7N��u*��G&�<N�vQ�q�G��eS���<J�Ue}f�B϶��Z�'�9��ød�z�d���:q�Q8�u���1yL3FMf�W�½l� @^nb�3�bK�O=#� ��G�Y�:�a�ic:�����,���^� �-8�፶ŀ"bv�]��(|K�B<��SkNM����5���s������N�A*X���I:}g�5��|2��ߛ�r�-	W�-H8�Ѷ�� Z���	%��+�yX�� �iۀ���&Rjf;����$��2Z������!,��ߚty9I�b�ؚ��a}�v�џ��7E�V����9χ�w~0pI"�b;mQ���0�p=�:��V>a����o(�{��	y=��*ئ-�����qƔ��"��d�����!R�z�TMgH`�"�B��ߕ�V>��p\�/��l׵��qR�[E}�و� n~�N��<֫Hϭ�b(t.�TX��?�9���̜ܓ���2Ȫ^��MV��n4($0q��Y	�+@��e��P����3�`c�2���V�:���we�Hۤ5����a�B���K��"i�(��~G�����+�)0�Y��T��A�r�zZZC�rO$D����^�׺��˹Dzp��=�^�W�>ߌ��>��d���r�^MVTtgS~I������~@3S�!{�;_�bV6p��E+�[�������	CL�ҝ�k�e�k/���z�wci-/��cs��RϷu�	E�W����+0,\��Z�Ǒ�U�Y]�~��z�iy�UI]��7�����d�o(ǚ��&����4C�ͩX�c�z�MR��VFb�1P�T@e��͚�9+p����B�w0�<�EEP;:��pvC2�\�@�r�]xh6Z��l�d�BKUE&E�+N�'���%�E�d�W�:5�d���_!��$�[��ś�	G�{�D]t��t��}�c���OPu�A�&�&�Tyح�|ec�]kF�Լޡ&e ����D>2�|�|�2.ܸɽ'�g��Fѩ�ӊ��v��GC<pcX��d� ʙ�:L��Q3{��A�sT��xD�X�/�6�}�XN	,B��.�7In,��(�M�`�>T9�,G�b�A��R�U�-���(N
�5������M������a4 ��`��z�d�2�,nX~�Jx���j%Ac4Y?7�nS��6���Q��Y���-x�U��Q�|[��9�Uj�����(!�_I���i��ZO�"��ITs�7���l-���83�WR����8�R�4x�zLy�����c�hyZX��M�v�1[O���ϕ� �uI~�+]7�\B���-�=��b�r��e��Z�o� 4a���A䡼�~�&��p_��:�8�{����V���p����\ٚ��s�'3n���(�?AtgOW�Y�Q�T/i�b�rI�b�*�@���l)���;�	�+RԤ�b�:?e�~��ÊK�l�7h#�:�h�� �"Z��/�ū�>o����㙈!�j)��̴;���\֨�v4��� �M�P��������P���߷��(�T��:vIz'_9=��J�;��Q��v��ˣ#>v� ׇ"	����7
`��~�������jU�|��gvr1�ar~��^�|\����t�\�6�uy��FzL�Fbgv��F��@Y
�X�Ӆ��%�-�/�M��1���47X(&���w�tλi�R�?᛿o�n��@���@�o��Y�R�������]�Rp�#����@y��AϚ�a8��(6Ӷ�����7���w��ιO�̍���?7�^|:u�{���fBw�5/"R���UVj���k�!�L"�x���?��ٟ�x�6�	)1VmwӁ���k Bg�ٓ\�Ro/�>���v++��4�5�P�EDe_)����M��e#���O�����S��	�Ji����ɳ��w��'Ԕq�p�FL&U�M�x@�=�{>ڝ�)�QD+w�x�XhO���u��ݧ�h��oz܉Ɠ	,#��sf%_/_l��RAX�7'{3�5�%�
�������6\�e<E��ȃ�5�� ��M�k��9�$l�*0�gh�UOf �/G�*ꁽ�UK��(}��@88�ˆ�O�����%��|�ǁl�T5�G��d�8v�~<s{�!�N��Qkm$`g;��˧c��3�C��^=�Xwe�p�
���=܊c*hi��Mh<d/��G�\̕��Zo�ȇ�����+7D"��@��V���a�(7��z�X��.O'�#G->yS��s��U��Ŷî'1����a����Q��e�+V���W���83�V��aq?l��$Lj�QT�b!Wv.'z���Q���g�d��O�i���,�N��R���{8��u��6͋�ݨ�:�97M�O9��O��$�$Q��Ű��.�!�M'�@� ��ɭO��z�ԭl����+J���S�%(�=�Y�������`�Y��L<`���x���'�x%JS�{v'*����>�Qz֗�8��:SL��m�ƽ��\�;�]ֲ�m|D(�2��b?*u�V��&���ne<�e]�gP/����'���Q;{���3�y)�����gH�~5�r
�����D�al`w�63�{Ħ�����ш�HS���0�B����Kc��	˷Lz��]���Z�Z׋��ih�'˟O�Nw�n2��ip�����L�l�3�GCBR#�-fl�I��ַ����a�/̓TT2 K�� $|#x,�a�/�?XO���\δ������F-���R~=��'#I��/*8��|��.��B�``�%�(N}G�+�Z��ģ�>������?��^�5�R�5592�*$����%�k1��ɍ���w����E�[\xna��0�&��X�rU;!�좐��`M���Mi�����"3i�"��k�80���Hf%�A�*���r3�b����I��?�>x�A�d��E:�Ou!���V�!�Y���H�@���&�3(�+/ 	��4]26P��<zS��z=��	J2,�o���TR*C�=�\;E���?����9�X���4�9�Q��׶QD68~?��y��*1|��ٿ<o��ϿJȯ:z�ÍN�	���,t��� ���`�`�y��:l��.�MR�����u-��^�)�j�'�v�wH�(�����b���B��W���mvc��߾̾��K��I�,�h+u=;����0�D�<f�Wa%�4�qե\�ggA34��Lo���<�����&0+�X����03cAO�X4�����56��|G�)6T��z+��uH��9���hc��X�����JV����H�=���@����zI�+\���%WEϿI���Rl.d��#4��)Fy�jq�RY��ϣ34{c���}��L��더e����G�rV6Q�3 ��	�C���������.��E���g�U��^����`8����g_s?��]��2x>�l�|�.��P�ɔ�4�[I�0�JEq�~�c��ຊ��]L2$�g!�����,Z2�~���iu��<$�k#[��U�������h��P6^*,�K�*��O�g	5`���zܨ@)\]����%�'[��&��u����'Qy+�aw=&1'��Wl�m�B��bT')XW�ZB[�;TX�������3yj���/��5��-���)�8�v����SH*�GS��^�������\�5����`���
Zzܗ���'}K{G�J^�9��<J�o��s���у���ؓh���sI�!z&^,'���y���u_T��P�2Rj�v���'��^0�)!^��dq�&��蔹>!	v��tظ�K��m	�PL�9�;׫a�/���ˠ��a4���G�U�V(�R���g!W�������5��4k��p?����Ea炒�EuR��`���\E�<�D{H��d8;����e��Hͥؖqĳ�%�����;Vsc�Y��U�hb^�0P0z��Wx��z����A�:內����镝cbjN/x��E���necx�{v�h�[�r.E��,�ht@�E��sD�𙮦�V�[���Y��-���M�5���ځa�[vhz5`;���S�v�j��?�����,�qdc���5���O���[�9oM��N,�p���[WQ5b���I�4�P����k����6�H7���T�P]JV���Ѝw��ȹ����v�<��_)��kP��O%ݓ#�X�W��qf��I�S>p����8KG*�ã�����^���_���V��~����jν�w�H	_�O�U�P���B��N���q�� ��A#�D����))DC���"h��8���3��7#����@�13OV��Lf�Ep6�D���eؔ�P=��<�Y�;��QKN��8���]�3�B�1̝�*J���M�l�U�V`�S׆\\c��c:ă�'uV�J:��P�� �ɔ�I�A/dUwK.��QW	2�l��}D*<���1��nh���JQg;_�t0���{�����BBP�W��R�����h5V]�}����hC��L%&)9W��?Yk/��s�
��X
���'�w�� +������$q���l����םg�E6u5��b,���T_������ Σ��}����-�3���E��y,D��8i���
�+>c��Q��ҿ���<O�>�7JZ�)g��׾uݓT�Vi�X���'�/����Ŗ�/�	�7���y��A���k7
�ZH���hK�$R.���R�&f��e��v�m#�+<���GZ�[��T@F���ʄK��$Y��m	������v�}�s� "�hx�G#��X�Ĵ9s�DFe�  Q��Rٗ���&j"N���둄贫h�rcׇ�RS8������Y$a�9��$=A��W6	j}���1�s�|�V��D�
Kn}6���?����Ŷ"�x��B7��h�����S��aP�pM�w�"թߏ?�G�ĕ�mz[������b=ɏ��v ���O�;����懫�����d�3�j�-i���ٵR�^���&k�Kխ_A�P�:L6ع˘ 1�����5b;���v˅`\\�)����S��w�~&�	�ZR+(�j�b�e���)4��<l��{���H.��tI��~sFvs��/�誰,7=R-wu�SO�A�LL���ڣ5��%ݮX�R�`+�G�����v�<KDrTH�oìP�2![��Y��i,�^�S��lOg��B;��r�`I����H$�*'��~7Հ�~Cw���(݅�D
+�2ݲB^3�~ZP������Yz�8,�$xr]E�ѥx��dB�#��@C�q����Y5���D�D�3a��|#��達�֔i2�-����,�����żOBhkLNm\�̹]q��d�0�	��䖂q���j�x�7_Nx7�[`}��	͙G�q�s�(�3��ݱ��sBz"�YՄUyA����f��:g�/���x����i�,����З��i$[[w�^�UP�|��-�"���?߰��<�^p�k�bT��`��q^4��OK�W���4�ƾ+�U�N:꠾���x���}�	lT�qN�j}�]x�2!�2����
y��G,�KG�P]�O�O7�cG9���x���%�=��Il����,|
�h{�a: (o�#��m>�VxڲM����U��\��
6��/D��6���%���h��C9�'b	���)R(i��%b���K'M�>9�)W�
�L�pwK>�h�L�X�,�"X"��Ƕ�f�@D����^�=ӥ���2@=�ҡ�J�4q�<�<��[��g���N��Q��������f��ZD�p�5R�1jjVe/]?nc�	��vz�x�b���(��4G`u>��*�tզ�׈������/�3���r4�!Q��gI��Ԁ��U�o��VT��ȌG.$q�Pw������Jhu���r�=d+�`+F0����@u �!����U\)�U:	ws�8s��XZf��)��b[.�	�86�9�m�e7����R�""#�!{�B���]��ٹ��)�^�G�sxƸ	�{�	q��B��y�n
r�5H���j�X>]f�V"�Sm�|v�V��h�K��'F@݁���R���`sy�B/�u�6�����H	�.��}��}����wH^+�5䭷y�F�}$`�~�5��l&W:�+f�m��n�� 4�>Y\��s�&L;�7h�H˴��N�sv���$�����_���:c�"WF���ħ���\���\/��O�F������bq�t?���EJ��i�#O$�F��Ec٭c�a�1	��J����L����.����t���9u����������t�a�n�̽�.��uu��F��n=���_FDL.�N�)�m�F�Ε�9q��p�'!�(O��`��s��e�� 7�<x^۷�k-h�5��1.+��	��@h��2y�
Z�e|�fzy�,&�*O]�}�yM�d��(���P���w��B@Į�"�����|�a����q��l)�D&���T����s�����d��cl�ۚ�abv�̧��*<��w��~PZ�����=3�3���d�����_4��྄V	z�m*�@4�*� �\�3� �u�F��!��u��G�{��W���'�S�P��-�7�o�c�{�ۣfz��ªT�Y ��ڠ���K�|�U�X��MbAՄ ��WrrbR<p��f��ׁ\�=UהĢq�c� K��g�*+��S����Q m{��b���!vYA�&"��]��y�Ԯ�r�=%	=�_[�n.C�T��#�a�K�Fʯ��-�TC;6�7�;2F�$�ƳY;mw�A��8�b{e�q��(MM�L]�;9c �iV��:�cy�RΤs)ZKS��� j���yO��x�I�aG�CڻK���h�<�L�?VĖ�G-��k#4(N�_/��Pp�:N�e�p�����sa�Ӏ*0�V`�!*q5�O�'f6T�h������%�ٻ�X�^�馤!,��0>{�կB��9vrL�I�c/;?��aC�{���8v~i�֨$+���*8~��EF�.�'�.9�;�!<�>MneV	�}����3�2�F[����z��Q�o�d��������+}G���&܎����6��x�6kظ�,+5������x^0*{e����<��5�1�3TD��~|-8����@<����S��~���kxU����&K\� Dn��q�dB�q����Y���0���nC�_7�2�L���n��$��u�gi]���:'�Eˍ��2�J4���tk���3�����Ѝ;w���P.IW���lC�3���6�$��뫖(K���PZ�E��:�� �������nq�����#;ψ�Hr d����c��oٔe�)������d��j���e�0X˷F�K�4��7^������ù+�9C�J���J����v��)
hN��Ux��wu;1^IK��&@�a�!���ZP�&��\A��;}]���&K'���v��o��٘�:����F o~,&���crS�����wf78�X=s���q5� ���E�
��HO�eJ��%��W�Ȅ�s�Rx�����z7��b��TWT�`rŉ�v���L��B�xǯ7m�p�IӞ�������[)p�0jkWaͪ2���RT�_Ϭ��͜UoΊ����l9ڵ����p�G)ϑH����Nw�*Y�J�'��aI����}:)�l�4�UP�-��)��&a���Ƿpƥ�m[v�@��&Vg���̜h� �Kh��k�cK�;�	%op!��,���������n��Y_�A1nl������ߔC"���j׊��e�Ct{��m�H��kg��W�s��+�I��)���J���%Np���=��c<�U	���򴛡����i�\7',�?F�R�tCz�!�i�/+��|v4-ŢL��c`ѯ�A��}�ܶ�GV1�?��G�q���b�_�?�����i�́��E���]IGW04 ���׍( �%w|
`�oN@0��k>�k�ɭ���Q�TX'C n=�(%_�&\���Tf8���t���/�Hz:�"-�Ҩ+Y�������t�dā+{��G�������_$�b����M�T�!7ǀs��3̓ٺ�g(#z0�B�WRI���)�a�w�'Zx�`(-W|���?8k7uH�(�Q�2�?2;2��dU�I���W�jô��'�X�l��� �UH3�*U���	�n� U���?�8�щ��o��;'������gv�خ<��TQy��-�^v�;���
�|�����5�R[�4��S%��7.��r�8�$1�����z�l�G�D�G�ڎ^hp�̎97K �3�D�f���h �U5�T!�e���mt S�On]@5^�n���Q�iYD7G�U�$���s�%�l¦- �C�=�k�
#� �ž��6��P��X��s|iMC�xq�#~�(��ؗ2�zhvs&�FZ��+�R~Y��*�~�p�N�kQ�4�F�G�؂�i���]�֊�����N�O��:�YM�m���(�K6Z�0�����p����ST�!r�ib�Uݾ�z�z\r辐{{�1ؿ�~���@/��gB���'� P{hV2V���#:�pP�l$�&2�ސ��hN�\��<� x���І~q��	T�vT�f��=�ނ�A�Go��H��լ< ���i���񖜠�{�>
�i�f����'=�uV���C��O��W�!����z(�Uy$\8��O�*�0����Pf�iZ���L>c~H�|��jws�	Y�m�K�]0H�i�ש)/����Lᒵ\�[���#�����3�6�B��}��ֱ��9'x/��RPo�uO��_�ɧ�<�^�3�W�!�z/w�0r�y��<���^�Rc=I�TQ\�2����C�&Rc�X<+�,3sN����;�ߒ*qtt�ne���c�@q�~x�/�R@���i�_��%�Z��My�ܲ?�}��ey7�Bg�jh�%�@�f�/�D�qn�Bc��a;.�}�s�ع��$���7�h]�f��7����th�s�@5
����n�Q� !��D|Γ��Y+����>���o$�C��`��y��H�.&KSZ۷|��R����ǃ*J�%��ٿ��r3���c�Sc_�!�� E/�X^Tq�����oRf!�Gm��q��kq�UR�E
{z���QyǄ��>@>���
�4.�&���;���_jnx`��^\�Ϭ��o#{���ZIR�)�*��D��I����kn]����1h����c�q����\�����$��FV��;��ow^�$�ٜ�*|(u�1��M͖n�!��IIrR«�N@�Ö�Qh�T�J��f��9Ik�r�v>��W�O
+:���&@>���a�Ɨbo%�֨t�����˘k���pٷ@����
v(h��HDV�2����b�)e�ٜ{� ��3���^�ą��0��6w6�>��$8F�&_o �ߕ��<����yFzbTM���4��y�7V$��_:�h�j��ԹϿ�`���Ш+���"�V� !]6[ly4c��!��91O`�s�h,�'쭉���}2|n8�;}%�q��܄
��t�r���7'H,~�f�2c2P��͛p�K�L��<ks�öI�H4Q�J@�O�/���Pj.����g�?��KU��}�Y�&�G/N�M�BB'Z>U� `����S7�WFtݰ/2���}��\D�͙�*G�A�IZw��s��x�ԯ�q�X"��a�D@blI��j����H�8)���1?"���a�`�jT��+չ���:zj��JԶ�(�,��u������]&�1�C^�xT:�Ʈ��<7�a��A�����'��B�3�ĺ~8�q�\OЫ'���ςmx�?C� �G�qI@�yZϫ<�k��o�&�s�'�x_��h�z��~8BZf�d�Q�ET7��Y�/�����e`O���{�������9z``ד3^	��M�A��G�u��RH�"�F�c:����M�����p� �5Y�77�Zǯ�5�,�2�/�2MՕ+�h������p��2�_�pN����`^f���?�R�N��m_S�F^��+�����b˔eY���}�1��>�`�}�puِ�؞�8�$U�A!��(%/��8�sg��PR� �[��U�R  ݄f+��@��{�IdUQ��i�������'#�F��0�����f����a8'�q�'�l��%\-�����)��Ϥܓ�t▖��K4 d����S�˸�㾸�v������Ͷ�](���K���]�6��L�+��f(�u����14g�o�=�Q��j�)05�/��s9�c��% x�R?�.Ї|-�m����H�����x��J�����"��@�t6:�*�j��|��a��9�@��|4�f����	B��֓�z���5�<��1�дM<I7H�>(-�7�8"�����~� �O�ډ )��D�Y)1���lz���VH��4�ZF�j��DM�+?�#aK!���x�8������?E���)�>��Wɠs����G��H�Y��[/
��$vB��@��雃n����g$�[�ls�{�� <YiQ��o�  ��r�YhQ��q��G�j�`B;bC<����Ϡc͑��K}�g��&Y���ta�)�]����V�.���μ<��2���r�y~O�Zr�U����3���Uǣ|\���&2E�:��&�Ns�p$RTHb���M�#Li��"��u�&2�aXF{�R><���v���<�67���,�1�4���i:7O�F��\�7)/�LU��zD�[�V �,o�����"�I�J{>!�x�)�N��
�X�:qɳ��#���t�@�^���m/\& @7��dS��bǪR�;Sz�'����->��NnVC�w�o':]�7k�Z��v*���R�������^��f���ԩ�s�o@��K�Sm%ND-�thV��^�K:��rgN��0c!�N#�]h���z�Ia���^��8�,�L��>m6u����u})����Sz^����x[��7ı��2+�"y��S<:#�M��Me|P���^���xV�r�Np�s��r�z/��)�&,��_a7'�-UVa+ܤ�	ȼ�-��kAh�vE`<��񕰸�z,0� "~�ɠ��/@���]�W$����J����r`@C�\;A��lk�<���.��⥆Q��u����Vg,�*������ws�[Id�˯�&���|�!��lD��2)(퇲u�Y�����j�6�ԋŁ%����L�ձ:"<��SL�1I*��uW壷�q�zyv��*�&��#��s���l�6�g�����R��R�I�p�iu��P��lj�ʞ���HU'5�����qL@���m9@d-�8e�+p(-��$9�m������}u[���ۻ��R���+!�a����J=�ooߥH�!_����6^�s!].�l����	,l�ldN3W�JY;���d����P��Ii�,��.=	F�B�ż���w�i9�J��VK՟��?�+�񂇿%��X��AH�����U9e_�hN��:+��h��9v��s���^�!�/V���~.��ѭ���g�M��ǵ�|�lg3o�l.Mk��Uj�x
��7�Ã2��r���s��D~=�~u���˓axU�4-�0@���#1���BT���c����a�i`����K�[�A�\^Әp�K߄��9��U���nn���X�̾���2�" 9�;�ݝ��2I������Mr�1 �0{N� r�����bXD�q�^cY����m3s&h�%��,b��f�5�������^I�m�C��^��	f
��5O;�ǟ�E���`r�
@�!~���Œ��@�i��e�9��s��GE
B�#�*�Y��y��F.��w���z�#���>WWTF0�N��L3&���VR��!kqO-K�5ݰ>ckvE�1܊�(�fם��2Dv,��pəم�w�рhp�r��>���>�� �s�g������;[>2w"������x����7����m�Y���
@"�_�{̘�@rU'�.߾4��!��		I!�y8��A ��3�&́M��,��������y㱲�5�����i>e�{�I'�  j��".YeE���g��4�$����J���1�(C��	l�S��p�x�麎�#���_[�2�`Bv"�ZM�a�T� .�Y��xe�3�i��>/��j"m���3z6��e��7��D�5���ZS��d?�$��(��i;&6H��c����f��"3P�+N�bA�2|W�N�t��,K��3�8���ZYZ�%��
�x%hM�N�l�ZF��/#Z]�F\��q��l~���z��A�س��Ý��$�Y3�5Ya��Q?�$���o�jHwZC��`�k��>�`�+"�RތRt�qh�R�{PO�]�@!�d���v�y!�v3�8pwoo�" ��t�O��^솫����R]\f"쎀�@c\��OSY?
�]9��niT�y�Z��T��҄�Wuj����4.�!�p����2ٍ�� 6̹G6X-6���Bʬ�nW�]^ �v:�bD����x�����PÎķ�x *�ҭ�v��}��m�1nX0�f���)�!G���S���6^�ufٔy�T_ꦻ(ޤb��g� á�R .���+%��K)*�O���%��v�_���;w�D'��_y'A�������䃚��}�$j�u�r�l��y(��V�1��5��a��~�j�A|��xXln�����n�Ȫ����޴5�Y���R���pA�S;1!�-�^Q�=#*�i��r#�� s�M��b2��?ܼ(����,�H�1~��X#��X7����K/�ī	$�YDG�St E'����¶\�o�����"��f����І�O�N�(�.v}�0��TO��
��0�lsz�4EP���������O�� ���랪F�W��M�o��()'Q��0����u<Ob�U�Y,��K/cdT�8P!ԅ��TZ�e��!�Ƌ��B�	/Y�</踘cJ�+f�������V��Q�:��e��� �s��a��N��#D�������FR�߰����zȌ7"�d.g+�ų?"=�o����e�^g���L
"*�:�]؞C
�$<)�k�@P��٧j������z���U����ۻB�:<�w#/�yG��l:܏x0V>�YJ|�:6<b,�_.۟\_I�^�����r��|�Z5]P���5`�1��8T8�;e엲�!��`}�S�j���*�}֬B�Ҋ�Y��+�Q���&�#mj	j%����wߑd�»Á���%q_���Z��uyh���b����ڭ�`8ح�ϓY��§���a�a�}m�0�����qs��)�����	8������jZKb+��1ZL�0h�`�Pa|��"&fnzw�+%ϑ-���
DSH��V����*�ua��[yހ߁�����K�̺a�����2-q��ߟ[1���z�Q�vqF��i�Ol�j��[y��haK�3<ܼi�M�O"�Bs_)'b�g~�p�l��mP��*ň ����7A��A��`��̮Ӭ�jB�)���żM1p�b���� �d�zM���}�"Ƿ��ɟ�O�����w��OV���Ń�XZ��:�z/~_m#L��a��V*d;�_���؀I�g����-@T~it6Ȧ+�֖�O��/�M=��%_��#3�Vmv�њa���M`E�_vą��3]x���[��vlT�E�.\��{Z��cʌ<��~�Q<��CCΖ�qf���7��&�BF㽊�!>��;[��&]�<乪o@`�,�� u�����HG�B��A:�8G$_:�}�IlC��`eA��q����o�*�����-�D"�}v�y�(��}�6w�
��b�*��)W�P%�ܸ*�E  %��� vg���
�*�N*���3��Bc�J"d�Uz:�����`u9�2b�ib(@�h��O�J�+���G���|6�}1�>�O��3�~ ���K�	@�v�?�&��F�$6�&߱w_��j��m���f��A�O�%y�:#���Z9�Z�����y 7r���`���_��|���3��/vLz�.�3��/L̤?: �j��Z*����k'B$�q��8vn���l~�w���\D	����'���,*��+c��@��VM�\�l���pEIʶ1<"^�*����7�n��r��>]��OhY:	�����<2�;j�k����'�n4����)��C�.�d`64W�2����&�@
�+�������w&�.�9!�"s��[zm���\ۆs�B�e=� 0&�y�+�t�����2��#a&�{-���65��j5�|��h^����y��,tDy�A��9��I|�e����s���⭸N$�r���#�ҲoXn@�Q��E������P�?�9��R�t-썉�T��,7�s7�n0Ĳb��ZN��iAn�?M?Y���>�C%��c��6 �80�;�k(��ӳ(d$l��Q��$���|[�5�Q�r7��~n�P��o^�d�J���>yq�^&��;� r�ݰf�T���|���Ts�g1���6v�J*|`D��k2�_&��R+�������f��3��q��J�sqD���!�!��YK���"���O���li����ǣ=���gm���^�W8����K7��YD�Hf��2�f8�X���[cǨ|>���]���h��}bO/��݃Yֹ���ݵ4B�`J�2�5�t�+�K�%��F������G��>ϖ��°+r�0E�;��#�h�Ɋ�E�����f�p�{-6Y��4�ۚ�SZ�[�q�&���"���O&I�]7�x�	�[�_Ya��͍���J��'����Ġ$�L�-&*.>�Q�%FB�k(���_`�������q�pwpkR�.�F�=�&zƞ���Db�UhD��f�9�|&f3Zh-H�)��,��-wd����c����\���r�u���[vBN�������2,{��J5D�&r�_��ߏ�Pʛͫ��kD�;�j"������N`_�:#�1i��H̹�����8�H��$�݆�K��h2`|e�� ��˄�n5L���w�5�y����¿��9��~B��9���"3U	<�j6+�?��B�2hzu���c%��Rp�\��z��z�_gΗ���_�x�γ�K���]���X��Q8�����<1~�����	_[�����c�DS{�S:�Z���MQ����I�빡�LH���y&�~���>�yǶ�d�Fɟ�/4����\4��A� �,��#_������<�@5E�mGY��~f-��S�FD���W��|.Qd����˭�8�ώ��p��Ko�FD�4�.+�� Ym�@���<�s'{��5�
�R�C�ܕ���R����*/I�q����2F�̓���)Om�ǗH$�BA	��`��N�ʆ��Y���$����ё���L��%��DUs�&s�QA��8N�ޒ�>z�sR��:0S���u��aS\-��׾�C"�{�`F���a+���	���%k�����_���b�3d%"F�e*5[1�Z�_��
����5���M�-�r�$���l5\�	���Ҫ�88�v�ke�QT�.���:�9hJ��<�g��#^l�$$;�m�lpB:͘�@�r�J�C���@��JcU_��.m���7�\����	4jOH$���Wi�2o��G�������7ٜ�?e�b���A�C"nxX�m9�i��KM�;�<����\�;�
�S���w��\�&�o���-�MJ;�V��V_|a}��H����ᐤh�UQzīM��3!(�d�ӕn�A�3i�]���}!�^��a��?[q�
��1Vg�2L{�a����{^��^��a��A.2����umh��.���c{��ԣ�y�T�őJi�5�DcJoAa�Ič�7�֢HC����:��m�|-&N3ڴ�nJr���+�.�Jd�a�7�;i]*�	r�Ce�3����;K��>z�S]�B�%{�B�9wZ��g���*�:xor�8�g��T?�������X�Oz�h[-9LG]l��yZ+�6�B��j��3�kj�y�9)�fI�Tm��X���c�$�^O�X���R8j�5J�z:����������p��K��x�Q��Ѡ^Q�C)���-X4,�~�'XÉ�ד�.�����!��4����9:�?�%&?���P�|ܪ���s�ZKI7r
�H����Y����"l�![72)�a+�{�˻u��"�!	��$�Oյ�ܸV�/�v�d�E[��YL=�<yTt/x�wżi�����`��\�15�`[e���J���Tg���xA'	��P56"w�b�3}�U��H+S>���k��&���;:1���u7�M҄��hcf
����_�.������0C�c���!.�j������$�F �	�*X3 �`:�\������B�."
�rLQ��tt�9p�����k���F��������͒x�κ_�r;���/��Պ�)r�t�}c<���C�]nM�Ji�w�U,\���D���Ɇ�и�Q��"6��x�/H�Ö�Ѷ�85�͌뜀�9�����c��$���yF}��q\�l����:��"�nBJ��x��HtC��6�/�٩�0�ܲ=#ԗS�Y#zM��Ô��,C��E0���枳�P�8#�.���kä�᜖�T���E�ŎE$y|�Z��W �T���\�w�]�*?�-�rq���`G�b̡?A/�/�lړ�a2�_w����҃���_�!c(��:+W��B�M[\�=��X�.�n��=���<�&L漘���(1��kW�^����J�_���_��v08i�֊�O�����ݹ��%`&b�W�w'd���'Ǭ#�p��"��oTY-Q=�DQGkYw��oA�Y&@\�EB��M��r8L��#>'�5�e��1yѰwx�,|#��Z�䝷�Y�*X�x�����)�im�����L-͞���w%'�i@�N?���s���ux�E��¹��շQ	��,�ʵ�=x�I�{�� ]<^�&<q�;��\���"��@.J�V���ERf{��·c��Y�n<$ֺ�#כe|���NM�.�Ͻ�6f��a�T�EY�zZ��~,nGk��-d4Z͢3�u=@ҟ��	q\�G�O�_{�^�K�6z@k��H���*����-���?�Sچ�oP`�M^�fĽ�'dO�:EA~���c�"����?2{�E�:��ck�i��W�ϫ	�i���&��L�e&���X�(,G�%~'��걼�!�.)�45Űy�3���p�CU���ļ�m�@QD\"��)����w��Q�mE*l<��f�'�9����S�����o�GK��!?h_љ�F@\fVu�Ѥ�yC���ɉ"����1B�+��1��a�I��ꔶY�yo&�����Fއ�pG���K���"�C<���A����� �:��Y�)��7��2��xd�~N�ݐ�����9�r1>�|�~~�H;����@��@˶p�-�_ss���Md���5��E�\pA\�H���*,l� Ws��w(�l�[ �����R(d�����'^��9*��(c�s�o�eu�E_K�O�5�F�Bo�%�\�X��H�H�3:{]OboN�)��vgT�у#"7���j>m�)����|���inɺl<����"���Kؚ�k6�8��)E�%���>2|��T�R���#�j��>�g��^���}���g��Yu�҂�� �55^ڙ�Zc
 �uvO�����N�;11��%���bi�`��u��Ы#�mn����RF5���H���a��+��1Q͒��n�z��JU+�?��$L���#�a�s��P�*)��XI���|��^�Eq�����u˂w��z��L����B��e���"Y�
KZ�R�;�Ʒ�o]�>���q���w3@z�S��߅�r�y�~S�켶��i�G�G:��*�����QG�4�8)����R��aYe�0M��F�]����}Iy�dJ�0���������y &��.�l�Ԯh�}L�?(���Pե������*���r�U��z���"{���y'���3C��������d!7Sh`��7��H�Q`��"��E _f�9�$����W�B�t^�����TI	'��F����\a)9�����.���w�Rמ�o��pJ�I9�߰�����Hf��k�qyU�gBt���ڵ����;ͧ��=��a�6z1�t�2��������~�$����V���&ēc�dIK�~p
��d��!Ϊ	C�FG�byI� j28��	F��Ƽ!�.�J����T��D��e�@�ק��(�����z�R�+Fd�V�:��ذ��t�*�O��n�l�G�������C�D���l��֮�u6�h�z��&FM��;+J㖨��
�Y��-�&����8V�7����g�kXท[f�8����3eZC�R�����>�C�F�eH}Z�J�B�_F�}�،���j2�(reОf�����3eW4�pѫ��lӵt�W��s��wZq�(�f;r �m<�7
Х�F6���0#r���T��D�����Q�!nW
���1iي�v�GItc[H�?Z}+�>�g�d�������z�S&��V�q(^C�l��w^�D�W�	e3�!9 
#X�ƄԶ�ڙr�>�_�%��� } ��>1?/M��Xp���$>�v�:i#@S\�1Z�>�[�~�	��$}C�e�d�v*�|d�e+������I��)]S�fcT�
�����-�GU.��SUPE�����ͅ�&� 
RO�]4�M���vڮ��i�=�,j�����aO�ŖϏ #"x���L���Ah�5��$����W{됮���A��q�a
�,�u��!7�� � s� h��s��IEk��A�$�?c�6X���ch�a;8>[Pi�@�j��1[(��VF���[{����w.�_�$\�>,��/��%	]=�����V�:#��&���k��CK�w�:$S%��}����߯|7q�2��$12�TCZq!�/Z���[܀�����(Z�~�¸�6L~�'�n�7L��[4�)�c��%-�?��~������d瓲�qxޓ�)�\*w��\3�b"j8d繌wN�ս�>Q*μfz�Lw|w������[e����lx��M��s-���iO��-���YklK��
v�Ez��e�=WLM�����u���_�.#7l��α��Il�R��㣚,�o�}�ևR{wR�I�/��Tj#��u���-��tk��IK\
�~p�%A�
�W^�@ ��I,T%�{7.g�.��]�^s��~ ��WHZ;�@=��L��1v@�D�g#��-?������ϳ����'eI��HSK
Rr�b�;�2� NH�F�9܌��fa�J;��'D�yu2vc�" ��� ��L'I���u�c-����W�|賝��a{3�9_�$nJ���R�q���n�m����$���٥R����!c�4��� �j�6<�+�{[�p2�lG,�������K�V���A10���e���o��Z���DBO̪6��\��L��>C�!� ��.d.$qI�g���k�D���8�5�%���\_�v�u'�
��dN��Ք��1`���~<MEx�J�|��==:
�h�{yc�V�L4 �'oK?~�4=ʸi��+��z�<�2�f:�/s���m�d�SO��&��M�ƕ�K���tYQ��+X��N�/xk����U��k�$Nu����$9��im�Q�.i'��'��®�&@DL�^��ib�?$=��9��-������%(��Èzչ�KL�(��MB�3�L1�"���8�l�̳���w��1u� ҈�~?$�v�������ǍB�k���V1i�t̞��1a����kq�Һ|��R�6���K=�2��<����.�0���	��I�+�`54� ���������;O� T"����۴W�b�>�m�g E -��]VY�_��d�Te�]t���iv쌙z�����9�w�5(u�jй��o����@�6��1�c�B���|��?j���I؄�y7p<y�>��`�3��'���2��K��"�D�d�Fp���ע���B�<G�/����d���8b��"/��9^�[V4�����gL������h<9�m�O�a����F���JDH��y��P���_�e(HU����.D:	y��o�a��}I��"�n�2�5��<ӻoHW��o���":�dٚ�����B*{r���dwv7�2���؋���ҟ5�#�tX���e~ؑ�w{h��u�z`	��xo#Wi:���<q.�U0��>X;�G(;�d��m�������as$��S�4�?G`_�T?]�oe�=���9y��Ã2��&�@򻹐��A�2�X�C��@�6���0<K��Ͼ�����y���?��6D��PSK��{���'^p"wǉ�E����Ū�ذ�4��	<����2��7�fpǭ b]Q�Z%%~�<���t��NƅJyZ}�T�����]ŷ�J�S>�\�������OE�����]D���� �w�KՄڮƵn���d�+��E�^�����u���$��;a��_k;c��LLQ/MR6,F�����!���F�O�,(���1�{;0��h�⹟�)�Η+�j|��b�T ����Է_D���C�m,�M�9I�(v��T�����:�D��n�{F�/'o��{��\= ��O�C��ټ��W��"p��Wۻ��A4�=5l�_��_�t '� ^L�w��)����
�4�ЃR�L�ޏ[]k!��R ��jRmm���k��5�]�ƃdӝ����E� �(Q;pa����9R� 5�~<9wW��"��O�*;�0J��aR.L\����X��}���c|���I��j���5�&pkZ���2���Ɗ��rɷ~��:�ى��6Զ�!6�wQ(A�;��%�H�W��Z^潧X��{Q?�	��v�-�/p��.L��'4����q�Y[?/{
ļ��Sx��<7�_���U�l�����r=�P�i�z�h_��I��a±R:hY̕F7�t��(�B�����z��
	49��ػ܎"��l��x�n�](�F�;[�P�q��buJG�/p�J�<֓�,��W��|A��S'qJ��;`عs_E�G��a�uV;�0RIfdYZ��@���؁U�ík�"
�%�{�3�� �K�bur!?��޲*�@v
	���=��	��>���V,���[R�_=�a�n�$���3�;��З�
�\�ga<e����k�s߀q5%S�]�M��\O&�����xſ�Xz�Y��] @����h9�R>�NםO��GD?q�<T(k�B]��I��mK]O�d�C
;m�������<�Pt�%<{gU����[p���c�����Ӟ����b5�7�j)�e�9,�R�bH�F�jF�쯓,��3!G5#��M8��9�Wv�OϲZ�C�^f�+]��ڏ�@mȿ��Q�d��,v;V��!/��1��N��[&b_��^�Ҝ�0���
��z��f��0lK�|h\t%-Y�_����B��|�Kc�D���D��5���ѯmÁ�`J�W�/�p��!c\���7"fm�-��L(v�5$j/؜��2@gY�f̋�����[�V���1�"e��;f\
���5uyK<	�}i���I�jH8���ԣ�Kp��Ƿ�#2���!�W��y��?�_c�tiTE�.�@�9�&�ɽ�M��-��e#K�b��<�[�_ �?�i��l���*׍R�<��H�99������lܠ�=�&��GД҄��	�k���l"�2�P��O;	 6�h��1�O�%
R�.:w�N?gg�ћ���✂s�W�O�,6gnQC$�_���fw6��$��޻�~��d���慣z�"��U�&WuU �&>�=�)��<� �����0���%�k FY8,�F)�$A�y�bN�?'z��	J�  <��$k�}MB���&|�<����	��S�`j��I�]Xa/b��"����GG,p�5�:zH�� =�&ٖ#����eR�Yaˣ���JB��+��ǣ�nġ��y�罩icSIH�C������qe=o�s�S
� �6Z�	�Y�q�+�ۇ��-P��כH^�M�����B)��L�%Sx�,���l
�M)�q_@�x]�_Y*�����>?�έ�9�5���[�@�+g���C������9�"(TY���`f�v>�)f���1O+�ʅ�ڮg�U�e�N��{/d��s�c쥈2�1C�U���m��	��̋�4��`�Օ> ��6Uh�pAI�ݥ�țU�/w���Tz���|�Y:��I���P���n�͔1Vyl	0���PM���NX����>)6fh�?Z˰��C��1�̶��ӡ��h��(/�`�ls��E�ڳ�A��:��'�cЇ�f��k�j<��v:?-�@9��ug��������"��	�oL.��� &�[3)���k��.�n�{���z�c�4i$���]��E��3�Fw���	;~�ƫ���1�N?���%TIA]����WY&��0��T�̊�R��Z�P�Q7����T��^�o�q�?�H9�كL���ۢ�b��;;�aj�W�-��D;Y৒�.yF%�1?F�u��%`'�YuoX�h��n
d��.�=��,<��F��k�Β��4�m�]�7��1�~dr�n)d������:�6�eW
�����HI&:���+�'��ٻ�%���¡���s�D�1.��*�N.x0i�c���a���`	rC���:�C@��C�P "��P*�>½G�J�8�hq�?~2��N��DվZR4KH�w��r��j���P�������B�σ��y�!t���Ԓi�����|WF8�,u��I����B�(?�u'}2�q��k��S�s�;HX��!��S��jP���D�}8ew�8����gϠ��)��k�Z�k4��Y���3�����SCB&
�0H(�M��S	�c=���d6f���:���p�!V��b��Mz�İ��@-�����(T7���ܹ/xT�P�S�a�<�ӱM�N�)X�J���БZMԒ�"�^�f�\)�q!�?3 �?����`�f�I��I����$� ����{n��&���+gʰ��q/�*\Vq�ᅚ���A9ے��G*6ܾtf4�.�5"��U�5V|� >�8��!��A�G�-������.��-��Tx)��g��I�"gR5	p��������X��Q�+KP7��C�	�\bF�i+�p�k`�g��Q�g["���҄?A��X�g�V� Uו��E�T��G> �E2��]x�b�M�z�?��T���|US�����iU�s�.s��2ܘ@�k��*�}�ڧ����V��_S+�d?4���D)�qk�%��r(��������N--�Of�?0�Am0�
k�%]�u��\c�K�4���{����x���Ȉ'�C��8�3�vb���{y�S��F'}*z1����>���yBV�7��$�	�T��k���3��x�t��N����¸˯Il���	���F����S�lҌ�������(�A�#|?_j��#li��F9-E\&�,�t*��>zL|ɦMm��:�;��7^�`h��0��7´׮+�@o$�&];T�ZJ7�_��Ժ�_c��w�&DXxU���?�ڛw���O�#��e��k­�4
�|L��]��?-�ԫ�Z���u#�U ��.N��}��b������&��q-޴�9U@��ɫ���p١E����hT�S(�\(�:�J�u��C̀=��7�;�)!��-;M�e���
���[ä_(re�?�����pL�(c�R��q5�e��T�J�E�-���(K�p!U�,���/��V����4��f��9{��f��y��eiSw2�g훬����=H�ª
BN�|�B���G�1i�J8�b�%/��^���c�<n�7}}�G���K@��HQ�6/��Y�Մ�-�:s�.�x�������W�dޞڃ;����:R��"��C�� MbA�_7l�=�׿�w� ��S?Vj����G� �r��~�����E�D��xm�o�cE�i�����I�r��Z����[���e���u����}& �MJ�Fy�_^fe��;'�h����	�iC;)`9h�d�hF$�h![E��Ru�Kr�fཋ���;��CS$��Ǆ�4ml�� ?z���z,?��S�����܇)(�؋��y�S+[�M��ܕ��D}#�k�V�
r엋�?�ü�Z����P��C:M�r�9vWܺ��ҊB��D��_��%��-â��33�����/��Ҵ���Dh�K�{�*�/1 � $Xs�;_���CR�_3����m�q��~�W��*��},d"�g�����#���7�GAf��umN`5e�X��W"�G��vѶ�vO�'�:�:��@�'�;x��.�@0���a�g���RR�ŭwK�>F@�M�ߔ��s��8��X2Q�i�	l�I�F��T�&',$!�����C��$/�i�s��K|�!A��ٚ��Ӭ�efrJ�	��7�uy?D{u$�����ə�وӚd3$¼�N�L��a(0����t����8�7���;ɶ�\a�Ibm�M�yNK��,��=�qv*/P ��
pK&.	�� �����X�ig��ق����7���d��`��	���e���m��D��N�6������qMq+��<�zc�K
;R����{Mt�.�9��9�8����Ϗe��O�����3PY����ᦿ�X�J������2��2�g�������.�*X���4�4����&��*�3]E]Ҳ������y74)?pE�,� �M�L�6�㵍��'t��9�#l���H/Po�����H�$�m9�����F�����H���\�����EhQ%�5h�����$�I��}N� �{�esW律��5�wU<��VR�1�����Z�-:E!�rX�1Ǫ>��xR������iI�D��N(3�֣`1�4�n*4���r���n9/��z`������e�t)y��!EB�?I�xsbY���E�*����3����E��b��̊u�� �R�m�7�_���k��Z���a)�')1����{����.X+De��eV��<g(6�w��p8B~ @�K�K�7'��+���:	M失�J<���/]&V��3Z������A1�6�}:���c��E��p��0�Z�Oƒ�?fŬӑG��ښ�?q9ܤt6�z�7�����.�koٻq��]���s�ږ7p��M\ mߨ��47��Q�?�3�0#��V(�"��tF`vRi��j{�h��'W�Y��jؔ�)|lx���j^����C�W��mp����U=�@�]W��z%7���-VM��w޾&��t?�I��&�j��-m,W����Y��Y��Jέ��!��6��~'�n���Lfۗ/��`�&�,/!���UE�'!�t�KB��
��ɦo敱��3�f y����VSL��4��~N]&�*Xש�XTiBJ���y�
�j=��3��NՎ'W���->�Giv76�/q�.�jA"R)�����T�;��܄��c�P/���|�?�p7N�JBAj3��F˓��Z�f?*H6�� �q_�Y^\��Q��a|ݭ���ib��r�B����C�m�F�n:E�ɧ��e&�L��"X��^��B�`Q��^lMz��[��������_�Ҝ>jx�s�Y1p�mI��S�k˷�d-ؕ��*�z�b#\����/T5s�p���X��i����۸n����(>�bI�K:G���9+{X1��֘�ǅƇ�>qa�X�]�6ܧ��5LE�����f�l"���E�j&���\b����e��I>j�zC��⦉S-n� $�M�ȇ��U��2H��-����i�� x��oq�_6؊?B�P��6�.��^��F�����W��H"+��r�$,H�7��L��s�9H��!7�h��lFTZ��T�.��(�j��C͜o�2�	��)��)�������:�oqPn��IE{c��t�j�%O�ǝ���_�G>��XY:��L��&l�Bjrw�/��j�Nb��ke�o�b���bg<ͺ������Q�0�^���Us���A�i��GG3k���k~��0�OH]��&�k�K��2CϮ�Pk�2�?���>�e�Le[�[�$ٖ&鎥+�O���i��_�o�:�q���|�9�P�נ�;E�KX/��{���Șn��o���:�����e �OUv��;�gSJ| 6�V�1�dO؎"���XΔ|"��lMo6э���kc	O��}�@9�[��WiPN�[��|�����s`��^�XiWYVj	�a𺒛�y�m���q��x9s���	�|St��I��)�-fAHOz��IK�r�{��+������ɉ�E3`iEQ4���1��@�Bik��l��He�_\{}�P+�zT,��H��Vq���PPC)��|��Ů���m�衯�g�0�5q�ܽe�9���:�>�R�#��N�"�X�.w��xL�x�i�م��S�5i� L�y܅�ʷ��4�SJ������/ ei;�~%��`F+�6q�����K��Y�����:(�Q����p�Oqg �y`�㧙�U5�᪔�&�� ��$�Q�[C����g`��D�����M \4�X�Q0�6�b��u���nY�ф�D�--a��t�2"�h�B������ay��{��K�F,�)W�k3�f��j}�A�n�b	�W��#��&D�J���E��}/@`N�V�dw�����\\��`��t��"�q�bܿjp�Ұ:��m:��2����zu/�dRް�b��7.�vN�MiKcQ��K4�l��6]:,l�����K6=����Į��a���=�����,���ua\c�n��,T~�l2��x���L"�"�%��DKnf}�~��I�����/:� �ྏe�j��n�S�v�����+\�kQ�3�����Fy�$��J��Țՙ���J��������Өy��U��~n�o��g�Q�yWxv G�I��M���@��h�q Y�wBl0vBAsZ\��7�c�/�$n���M�c��YϸN;J�]���r��t�������})��zD���_�0��}B,�ɂ+�0ZG��b����Y|d�0��v%���Eo����;�אi��u�x�߈�^-�6;�f�P�A�@8 ͼ-���I�#Mv=<�b:x�l#dj������4p勣X�M�7˫�O^��'�鑻�A¯nE�VJ=`��a����/f�:�qh�3�rz���u�g~9f�b���� ��[�%��NM؟���	N���\e�L�ߛ�^ YLC_�Zԛ8'��nVNC�սK�Hw�Y�[�����sĜ~����L��:@�D"Lo'��ۚX�+Uo���B�V�)t�0���|�=.�DR�p�U�q�rɗ���^m*�g�`g���������s/2.aT{�X��-�ɥQ"�KE�پ��9��P!J�5���v�Tцψ��o{�.,A�!,�[x���T1?���KV�v�#R��{^����6���i���P�3����Ƌ+�A���Q�)o�;�#8�|}=S��ׄ_�e��CJ�#���@�$⻮�<n.,�/��^,�rU;��qt���D�Wa��sX�4U�Y�w���4�d�XDՂ�v)k��KI�, M�����!��>�EM��P~���H7�����+O��� S���&ew�5���r1���}�ٕF��p����ݏ�I"ՠ��j��d�{Gm북c���N�Oi�B�D9%��y^��U�"ٲ���*�k�oa�F`���-���IT��U�����e����C��gih8�2W�`�,o�DA盯�'K��X*��ڡTx��Z��q��O���d��d<X��Hn�������J�����Jif,H�C��`��M�� �CgD�1�[�Xӆ��:�it&+���L���#W+�&2M2gO��M"H�S��E?�np�R8/�3��#5��fa6��z�Xu�Qh/�	�"�BGA�[]�1Mt�>(����r:oi����+m�k��˭�ZW�X�� �>K��.�)�Rn���T[��9A��-ż�WjR�*�_�	���]��GeȤ�D��·����	���ڃ��u>�&�H�g1$��aM��x�(�4b�t�:ԻI>�Y�~��<!t��������m0��C�l���w��9�o����vQ��tώ+������T$~��:��S75�ʆ!��Ϯ5�CJ�Ҽ����/��h���"jĳ�M�[�����Q�kw��S݉Q�J�1}��ɮf.�۠NBKz��� �����sDW+�c���"1e�m�L�>�,�,��>����FƪiEGޣkէ�!���1�C����=)�2�Y��K`�jg`�m)`��4G� �|�CP3�St$Fc���3j�Gn��XwF�*�<cu]�v�I�[�xz� �`���0~t���R�s���3S��/2o�S�]�%�������Bö�[�^S�6��x�{P�pL#M|'ƯZ��JT�M=�	���Cd��P'����3e]�T��8L����p���j���8b"vr�B��R�Η��p3@�zj��������h�O�g���],p�g^3^U�S���%��E�{z�V��0��8��N(���K��M�>�Ҁ������uA�W��Ɨo���8%����]���q��oP$�Q�&�Y`�[����خ?�n��ŷ)�i�Ns��+K]�V�k�P-ϴ�(
�]`\S^����������F��,������9�G����j_>����M�͂�v�>^�����#�ۋ��R�=j��
���W<�C��s�N%ď�j�`�)�>*��ܩKN�^s��1�����,�4�	����:sLv!���4�ة����Ѩ��OD'-a���\������cps�lo��0.�MC����N6@������?I�G�R&�G�k��A��y�x�(�f���s����cі��Gv���<��Ek�[6��������caͨ���u��P��� �-����0K�F����{B73��Z��hR�H��C#vd�j�S��sja�P�5�`�9A-q�E ��k�b-|B�Υ�{L?�O�����ʆ���7�R�;��U���c�����#��������!��N����k�}ꅒ��G����t���	�V���NER��-
�7�t;l%������vp�0�(��t�� VŨ�G$O�����0
��Xq��?ad���ƣ�a��~$#�&�Lߜ˝�@D����=9v����9�b��=%�'��ކ��m������ye|��:�?�����`�=%��+W>-�]�0��r���@�>�I@T��O�~qG���rj�nR0t�
<+<`vE���R��+�B�a��{�0GW����"9M��S#�(u6��.?+{L3Z#��OR�*�Z�!TYjn9���(���r6�B,�8�:����n���65XР�RD2����r�+�,P?��$92�v��I��3.?��	b(�N%������z�+{�+�<�
��y�r��H����ᒽ�^�R~P��
�a3��ϛ��^aͩ�#����;��z�٨q��3����1�E����fպ�o7
鶑Y�
}�y>�7js��֊��'lp2�%���و24Z$p�\%�Ofv� �������&<�s��cT}��)��sJ�?]����U����~��g7?��~40㓚-~f}KO#��,��i���@a95����C���]�uR�F7��
?�N����4��L���b����^��c�7?�S2����(!'�bY���K��w��v��u��NLVHp��Yj��7yp����+���S��E�*��~���V��ŘRj��X�ܗ4G�~��0����Q�3#����ѶP}~&�D���ݨ��ۙ6���e^c��R�Lv�^l��9J��Q��8 ��ah({�*��O�P�I��^�͎�Α��Ł�"ؔkL����"xj<�YGQ��(��T(s�$aƥ�9��,
���cP�$�^�]BK���SyO���׵��]Ƙ�H��5�v��v�4�g^�n�x�+��)&.���P�<��Q��w�*<CM�M���4;-��)0J�[�Ѥ��\�XC�:(��+�Hѥ��@|M�Km6x"�@�U�8ܧ7�}C��pG����� F$��6�#��OB�X��4�FL!��%��_�r��PV�X��e����5�\�}���	%����N������n�	=�RIy]H�B����̘K�pwcj�L����YY�$	�क़{@A~�}pϢ�5�.3|��l,*����V-Z*�]٬��\���G�C{`y�Z0�}���]�i��"I�'Hw�	��J��������"�
[@��A��6V� ��GRm7hp`��7��G�b9 @�/�)���{��*����܄x�>�a�$��� ������ԣO&B4UG��3�P7Z���R���K��Yf����p6�M�,23�[s����x�Hl¶I�ו��h�O�w�جM�O;C]8ҁ��#D�.�K �TX�rJ�<�_������4��Ҿa��	Ce���
�B,���-jԔ|.��Y���ن�{��~��@nٮ�?�����0j�z;���w�,��eq{oJ�O�A�̎сۗ��p��H0!��~�x,�сR�ZHp�^�����ʋ�Œp W�v�o�^C��V3G�Ҫew��EV�CO�ۧN�б߷�r���ن@�f����t�Ib�2כ%���q@�D}G꒨Y�2�عp h��;�Y��f���@]xM[C�e����9�5�OTڝE&P���
��ҮO�%��ŏ|a"Q��f%�Z�9��3�+2��L �*b��֬�=x_~�,ZL�E�v��W�n�K.���ّ9�-�����>
�5w��>�s(J����u��d�0��wŻ�P&hÒ3'f&�1��@	�&����o��$�(��(x�DN�����g�dE~5�,^Zh�A�\~�h�t+���zԻ�6�/�=� �����7z�W_����ZH��f�����|�fmf	_@��Ƿ'J} �*�u��̜����ΐ쾢ű�c�=�"a�@HIA�KX�cA�i)іqkH9#�а�H��Z1����/ϐ06I0~8E�M2�nr�/��ؠA��rV0{�V|cS\����pl���":��Ij�KI�2��D���,��K����S�ɮ��+���8w�2�������__�1֒��v����TO6��*��A��[�cC%����'H+1�l�U;��D���pd\�Z�L�Ҹ�<p�_ɷܺ�9�1�"+���.�Okڍa҉��F?X���غ��<�p91��۽��Հ��y��38zS�&\w��1CSޏ��)C�Х�|��t�Ή>LI{.䱰�:"�������j��X���=�T����"T>��;E��\�.[ƒ���:�V��=*����������o_�%�`wyE�L���� ��M?U�3V�lj� �]�XK��$��G�:�oX&�D���b�(��z| �ה2�-^>ѸC07�������s+����� 2�a��v�&��}�۟9�$H��JHp{O���R� �2P&�K�_3��U{H�I�_ħ���ĳ�Bn��'O/��ш,���ذ�$P�k��}y�q(��p�������2j~�J��{�30:2hK;:�%�9!�>�Lh�Wi�b�����Y9�ZI7 �j�q	m��NE�m��WX��w+�0Y����B�������v�f~����� ����s<�Le�L�^T��,�[�G���uw�
��4�
�kB+���ȵ�_2�bCvCiQ�t�g���=�l[U���Rj�������wr3��=s�eR�um������]`7@�R�l�>�dZ�A�*$�1�^�ܕ݇j�iiۆX����>��������~$Ty������ڽ��kg��_�B�߱<}�?�o�����S�Opz��w!�l�d�W�y}�:��x{��9:��4�)z�ʹw�qa�P�Xop�I�'�����K�D��W;�XK�]� {���DC!�
��ճ�q�'����]�6Y�~%��F��}4�3b�RE�k�[}qQE{�IA�_zk�~�mz�+ �c�ی&�4�`�����$B�r-?h�Y`Sδ~��a� 6���v.9���։ފ#2�\�e��1�ĒX��D�h���WNFE4��aH�__��+N�v�Z4�)���JZ{�U���ϝ�Dn�e?�F���}��5y�E�[LkBV�oP=ֺD'��_6	Y���]��{�f@n�O�,��0��J�W�Z��;=�f�����A�Gl��`d
�Eu@f��X�&�o>��	
��-�����X;��UA���V@�y�^]��{��e��R����As��OT�qҊN�v�]9M��_Kg^)���H��:�3�߅h�z�EQ0k='�Cb������bݓ�n�˄Xa��'���+N���Hr�r�E _�K�gG����t�h�~`�����$b6�i�|���9N
2DJkX؋���6Y�,/l��q��c���>3A���74n}C�:!I�~�U�>���}�`�� ��^�s�X��k�:�0������jc����QW/ʼפu�BQb����?c>������(_@A�����ce������M��G��������CG�Q�o�XZ�S�s��~{\�n�wJ�!�Yy�H,��ٗqA���b
������K�/�w��9L�t�K��jYr dȰ��S���;���K2��,�M��b5� >!�^�
K�5lL*���'B����@�� ��Gƾ(�ʿ��6\`�AK��F������P��I��[š���[�R���C�|�U�N.�Y���t޾�����~��0場z�B�ڎ^��%	=��Y|�[�uZ�ń�.)r��:��9;���=�R��\��gİa��v�1�#�8Q�� w�s��~]��P�K�T�,�Mx�+��;ߐi�9X|j�W��ףW>�ę����wc���/���TQ����u�<�*���#�WdF#ɟ�8<����zb�ǀG�W(v�e,m���5��h4\šC^���4}8\M�yϤ�#��O��� �������1J����0����:�m u\�1�"7�������>I���wyrk�)t��i��}_%�Pr����|� (T��
�B��O�p�B��t�YԲھ����հ9�?��]�9cw�:�������5)�j�iU� �Zh;5��8��j�\I��&�ԃ,�����k&��7KJ�ժY*��2�քH泙���ێQ;Y�'Sֈ��Њ@b��t²C��H���Ap���� ���#���Q�H±�R��Yf�C�b�t��J�;����.U�>�=L<�
��x�F�S����3A����GX�e o'K ��-0!���9�^�I�� �����ϋ"���;��&o�L� �DvT>��z�g�$���/���@�-��P�+����G).��k�a��tYQD6�D鿗���]O�	q�'���ISf����|�u�	���+�������~�����U�b_��g��r3�7DBK�^=V��	�lmt�����a��=�9ވ�v >�`��w�)<JPc��6�`�?�8�;]6&�\b�B�F�E���p�7�߿ Y!o���?�x|�W�A����s�%�/�E�<��Ri���Q�j����� ������z�,�u6��i\f��D��`�+��U��y]l��lk5fR�l����R�؇2Z�?��R�)��Fe�Y���"a� ��x��ҧ�O;�`T��r6��Q�0h}���!�H��D�'�2�2������K轤] ����Ռ{;�D��gd�H=P"�?��y����'H�0���Đ	�~f��n�@
�B�y��J�@�$|�qG��3�k}fJ�� 
N4 �"f�,�&e����b��ӡ���L�ǫfY�M���_�o��gNS���%�Xߓy��`�}
���>��T�+gK[ḯ��Z��V���lL�߁j�����Mw�@X��\l]ś�5�T���h��}�G��x�Ir�\���6l[;V��+���S=r�ŕ�o��V���L�@��b{����c	OT"�}�m{z�L��rչ�gT�134Imn2�����r:���Zw��g����]<Sψ��ͪ��S_Θ8Ozڢ"�S���������u�[���f�AR	p�/�ݑ�Vܰ�"N�u�}.��(�ҧ�G�
5u���V�sb��'�%�.��*L�Н�&U�op�.ͨ�A��}a��`�X�U3��29�0>�7��j�9��
�=��������8����QrLS�����<����HTy��z����w�m��O����vʹq!� ��Ѫ���Ҫ��XCz�}Hb��3����XLNߙ_	Pb�N�}�zZik�M|�2ϓ:VdV�>�m�Y�ww��"O�0䤿�[)�ГKl���gcv|�$W�p�j4)8$�	�����,�Re�wӺ�3�R����V먵���a��8�*���P�'k~K�|_���^?B�{?��?�;������>��
;�����G���[�c�����9~�L?cxۋ?��ݍ�s�u�i��Dd6��P��4��t��[G����Πgdg�aI��1��:t�%g��]�RЋ��'���H]���J�"ܩ�*D:�a|��(�gLP����bO쳝���t6*�o_B�IX`��vA;�b+��a�#��0)/R�r�����]7 ��tq�=_#��`���/m��3F��nZ�y��rW�)޿|�XR�z��<�d���%�ס(��t�,�{8���9S�P�R6@S��gyK.en
��H������^�1�/�ajNޞIC˱l;t���۽�[Mpq�#�)�<4�=��P6� ή����^�ݡ���y�̭bkO�_ ���S���Oa8w�yJu��O���:��IR��{�W"&��\s� �N��m;Tě{��\Fehh�2[?�u+�aSJR\���(}E�We��J"(�M�p"��?ߎ���>��$!e����A�U�+<�=eg/=ŔE��w�p!��w��u�	�x��/"�s�Ψn[�U�絤T�ϖ�q�S,�߀?A2���T�W���Ü2Vǯ�y����ڙk`�c��U���O��t �.�n`�����N�b���P�\W���C��j�T	���F��d�����;�qG�U�̻����*�������V�NI)���'6��C41�r���� Hk"D�ȋ��ZО�W�����
�����Isև{�˨���="E��V����A���t$���zY�>���/@�2H�kD�L�U���s�P�,��ǈ����V�@����� ;�5<ɽ%���F�m~�ũg��=¶�D?��]���7!C���!�Ob��7�AB#%�!�|�\%R�[:�P��گ��81>���{�>�3v�����G��&����
���}�(�E��8G�F]Fw�^k�pcr6ˇ� ��&�p����W���u��wT_�^�؋1֒%y�pZ��(e��Fy8t�/,dN�q�j�Vhl�1��a:�Zr�Pf������)��;�J.<�_,��G�~���T����R+"AaG��m����E?��ܐp�Y�<l�	��Q��ǲG���и)��s�Z��v1����XW��&
�\۳���`[ֳ��<H�g�B�H�������`�%�`G,/Z�wd��8�e
R�3N@��)Gx��b�'o7Ф���o�Д������j�-v�ذ�WZX���~��S��[K�J�F �g���*0|�@�R�b���`y��x��@ݳ�He������Ao��V�lu	{i÷є�܏�R��8��*�]h!�lq)���9Ħ#��:����t	�]��ʧ��묠uB_��8os/,���
c�����%"掸^�vEYQ��I�L��L�?~�a>�A"��|��7gHb��,�`��7Nd9��*�K�p�"vo��0���>��u��8���L�H�߆�1���K�;	I��������e+`ʖ�v��`:�����G�"����NbO%��� �.B��)�;Q������`-��5��!ԑ m��(q�^D1/��KZ�,��6�]W�\﨨�PM�QNM��)�2;�x�IE����Ž��6�[a#���kng*XT��Y%+<\w��G՗�˂��}�m�.��lB�Ze�ky���/��ǽ��E/���k��c\�J���QaoVz�Sb��p���������Ժ	�,��HY\2T�>��W3	����S�e���)�.�-���:?�������JF;0�*�E�e���I%�G|�gvb3�L���m@.Ƈ�x!Z֔m@���V��_�#����|�2���<o�����4g0�>
vt
�8ϣjt�Ygm�'��󠉉F�c�9�
��GT��>���dhp"�^;�(B�@�Y;V��ɄB\�I��+0l�-�3��4������rO�n�����+0���'��t�8=��A�K�+��n�T���	�ŭ�,����)��6��2PU81$ra�Kp��d����\�V���C>�}g� �2jO�zmɛ���@ =�Y,�P��Lb���
��_�ǆ��1��`.�������:p��}��~���f�d��^�'��t���n4O�"�Y�x��~*~B����E�{�/��kj�����bѽ����x܃��
`�cjۧ�xLEc��K�?Jn��}�����^zC~%���N��hU�r*����?7��q�N�5��q��)��
h��1�2�=��6��Cl}HŲ~��^%�Ŋ�=����~{e��zU�o�ը����O�ʁ��8Q9��3����tP������e�~���L�Ng̦��)�Y�������T�'J���mN�es�'k��|eu,Y����K�r��:�cb��9}7t�ß�N"<���v�e�y��� m�?4`��3vC�#��F��v�idi;n��Dsׂ�R���|٦l.)��r(i����u$��^9O-�L��#�\
�<3�n�A�)�R�t��񝴻�1���
k�'c]cP�q�M���49�>��B��#;��s�K���[��V�*��F���<��ݪ��.)�o:��gVX��#����=j:��g�v%�l�A��%p�����N��|�#��G�8�<�Yaiw./d_�g����Щ%(��,���y3#��Xa�p?��Y�:E��o���3gU��r.M�Reͱ/ ��'��iqs����ǫc�����a$�hhJ�短Q�tőک���F�]�d�]�;0VqЮ������l�ݤ���[;��k"m���þ�Q[%�����S��L`n��TL%Ko�6e[�������c/�s��6��bA�w�^��EH�6a�e���t�\.r�*���(�3~��[�dp���	����߽�p�	�#7��^U�K����-56���Al��or`k��OXA׭�� �>!'����5�h���傳�� ��gS��dE�n�o�
K�XL������8)�&[P��_v�b$���!�DjM�J��#�<�$fI�Q��80x	/����`��w��=�%r}���'E�����#�����JH�&��QO���NT\�,�����/8��`��!�u#�o�j�����y��}[r�W��[���ڤ(��@ۨ2�����qJx`�΀(S�]+u� P�t�;g�%N�1$��oH}0G-���Yl[�L�<h��n�m�c���B�P�(?���P5���^���+�'����`�0Il���C�B����������4&2�K�;�FhȇՋ��-�9()	�tA\���:hhș,�tߢ�%���Q[&�V+0�,����S��
�4��@�n��b�ӭyܚD�{�f��a[��S���ˈ^@��YٳP��[I��D��kAd���/�|W�SB8���8x�=1IL��劭���N��jv��(�2��,+�&�QMbR�_W]�S�Q���+��o�������������D�&鯡���z.@��98���v���j��{Ϭ�f�ˍ�K��%����K�z�KqT���zP��\2��n0X���w�o��FQD��e��:6�Y�nXL�l�c���L��h���Oc@:7����J���~$y�"��/炈�^^�������(������\�-�G���˅�"5 A.� {�r�8"/	�9.J^>!�M�:E��n�(k%!*;�Z��ʃ%�6	�m��i=55t�׺�z7��3XE�փeȈcn՜A�q?e9:I0ָ-(�{*��_/��|���o��2;������ub���F85kB�İvrv9��'������"�P��_��������7���o�mկ]�S�.:����G��q+D������7��w�a`_3ߖ������^	����l�eD��s_3r�{�!p"�S(vN׋/��J��0�e/	��Ȓ^̛�t�MRƌrW��@w�#;�%=h`6~�����B/��˿:U0�ijS��rP�;�O��k��|z��Ӱ�Ҝ9RX���5v����/}��i���^|*�������SL߅PB�,4Ld���5&v�:��U�W��:5k� +�!�[$˼���T�^��[�D�-L���`$b����83�(-yL+/yҍt��yК2n:H���K�K�t�l�B�3A��*�����P�=7��Sg�F�^0U9Kt�{|Ղ�<G.�� ��.��k�{P���ڭ�?�%��9����-�׷�+X�֙�Ga���!�pL\�����g���pp���!�V����^�ΥI9�y�c��-�K���y*�]�z���T���L�}|��N�A8Y'F�����./����VғJ5��gлt��x[�K:xiq_#>���o;���@@A�ǥ��@��.�J���2�,|�v�2�Uc�U(O[�ֽ<f�����*f�i;f�ʤ����ſ�~�mbf�[Ǿ� p3%.	~�qv$-�1�|�y(rۈ�6*R��6w�t���5���~�`?WJ�4�䚝!�����������ٙs��f�,�zi�mc}W�}�6�:7���Ƙ�����f��Í���[0l�����;-�ǫ�����nT����iu�l 7�5�E���BG�B� 5��BH�;Q$�h�d �K���Կ�{�?�� @�r�1�/Uy�m�e��v�H��������m��_����J�Z�4Gư��1�P07�����	�.��c{&��4Y���	+Kn�u�㮣�ބ�� �ʥ?wр�N?�h�O<� �:�*��p�~�=��V��hl��s�������d���*-�	�l�M�f c�i�/��vt�J�����E��m�$�D��
q�S��p�k���V[��y��J��y=~���l&~�6��)r���>���ؾ��;1��rb+��R�66K�EX1Hc�]���lyV����E���}�b�o�m���p)n�����aA���f�WSD1f��;�L>z7�'=�D���L�f�c+���|�0z���|o�L��ɘ!K�~��k8] �XDTr6��*yVCib��քp�g�(r+�΍�O�0|o��q��=S�Q��W����+�]�����#N�e�H�m��d�:n��ݎ�������`�9܄.�~u��Q�/��I��٥���{��\�B�����X}� ;m�l�Y�h�#M���$1»���d٬�hd�몷�F�&Ä�#��]	⮩���M��ː�ښ��O鬧����4`c0`Ib�����ǉɅ�%��+H��5RPU�B�i�Y$r��!��E�N*5�L��'��<����u�Ǎ ��]��0����5�I�]�t?��G��ކLh�+�]��^/���Mٚ�Lz��z��0%%�x�j�T�Q�̀+�� �Z����������a��Q&=h��;��q�ݣB�~�- ]�Lv����ՠ�����
Y�=���"ړ�w���@z�D{~��Y����EJ Nƛ�#���o��t�������^GLZL�N�1��Ζ4+?� C�M���.p<�,�l��L) Wc���\g,�Cqn_~���;a�%�y�2�7 �ɶ��� 9���д(N9����=x����ҷ;t�n]v�O��#"f/����
�D�B�i��&ɕWAeRZ�o�<�� F6���14�`1p!y���啾
G+٠�_|�(����>��oǹi��kJBP�ϊA����H[����8$X��/��%Ze�9��PT��C+� �y��e?����5�a�z�K;���O���w*��ZmG������,�zDr5��OKtm9��G���k-��h6��������!?�Lpڛ.עu��M��T��Z��9���[���������u���h��:�f~l;?j��m)bvu������g�*A*��*�_U��9��~t�"V���!�0M�k��@d�@1�m�L�"���4K}�P
�����_�lg���;�a��Sa�f�e�-�U5�-�0E]�â�S���֧��{P�
�R�yp]o����{�b@�����n6UV���K5|^01���ֿ���9KR2Ђ��/��b��8#��`��voK9s�G��k� �n��c��z  ���J��w+1Ʈ5�"�Mk�c�G��W�b�Zu���o0mf����>]�#�a�öR�$��K��*K�c�ˍ��p�t־3 f����T,ڏ�1�#�����u�C*�ɾM���Ү�P�B�9��ǔ��W����]����?�MXI�^˜FS�$��ߏZ��4�'Xu��@�H���+�w1u%8s�!f���b\>��"7j�[��	�sIEX�=v*.���,`?L���N'Z�\�����lX�$k2�I����0��7ެwP�;
tU�#$�92���_��v���������$�Q#qEr\6�D���~��X�� �?�m*�����}����%����ڕV-a�ګ��ߜ�J=�Y�?Nݩ������m�r:��	����y�Tge�T�w��_��SN�Y�1}K���v�))�+h� �[�:fr�~l�3ΦI�*�Esޣ���������(y�.����*\7���k#���f��YtÊp�tX� #�N*�I�J���Vf�TR1�U=�F��#>k�"��S�>����g@�����=�ބ�鲂�W=�f�uo��pTMO��
��l�>_>��G�g�����s'!��O3�vp����v�&|�}�3	4�H���|���(�Y�]'�ݜ�3��Մ���C������k�����q��#���{�n�c4U�Ҍ�=GD� �"�lN �h�y(+��ƭ� �;_�/ɥ5Op���\>��2������&^�[x�p���9�"A%U������%�@�M������RF���wI2ͱ�IΊAi�*�zj��[��X���Y�-��@�!˔ςPk�uy;��kb�'@,����ϤM�[$-�+��D��� űMZ[��,οvb��X�36T��J�. s{U�~#H�[�Dy!�Z�����|����ǃ�o[��~Y�wl����yy�=1[�C���(f�%���n:O�Z��0K�;�]����7_�-E�hI���)Y1΁�\=	4��@m��M#��T���4%��v�1p��-�����
I�19}b?��t7Dz<����H1��mټ��֥X?��wsp%)�AUn0�,L3HxrǱ*rc4�/���s�{�Z�����˽l[uezTA��l�m�6���]�pEy�8"$&G�C���B�	 LA㦩[~��~����|��z�ؿ,O��c�Ӳ��?
�(p�?
����P8�e�7P��ڰ�F+�e���Iݔ�8��O�B�dn[O���D
 ���
��� �h���;��.�.S8	1w�Zh���R_����{qI�HEt�;�&S�Ԑ��8��;u�1�L���eB7,�x�	@�g"{���X� ��SQ�`\���Ըm�uWuT��8 \�=7��}P��O����1d�_�������_6��]��X��s�E�����ɏ�_ 8ie��@}����%x��I��`=�Ż�����jv��ː��^��&-���!���~�2�^Ue��i����%�<��g���OV��*��&Q�u��3�=]��$��5���Z՟����U��Cr�B�(y+!�d �c:�J�B���,�VZ$�"y�4�2��Lox|۽�g�o�GnF�b���������q��'��v�q��dܕs�r���o����vE��\��!I��#���!T�@A�Ϩ�m1�������I�e���	i�/tˬu1�l	����\[�S�ּ]Is�U-�i��s��5LO�s�]������V;�.AU�g����"sV��>0@}�i�fn�r��#�M�͂��K���f��	��݀�A��c�A���뻠VBe��c����G�$��E3����@d<㝈�Z!��4o����7��}�NmH��t'��C��X��H7��\ �Sgm�ɽ�;��9U�H��VG�3!'�:<��st��_��T�Ǆ�ݶ���6@c�c]$�n?�PƮ+{����F�zI�N�"������cf��ҕ�Z���Jɞ�Q�f��8��M�>�y�`Bt����A6!����a>5����%��HVxA:�A�`rra����Tl��J�g˗I�t|:|�D	���
�7i-g�gu,:0�F�y�.���d���H�[q9�!��M�pS;F����ÎU�-&$|I
FH���XI6��<���Š������1hխ�	�KĶ��V\'&��̃pU#��� ��H;l���M��4�Y�e���΀��9�H0Qͧ�@h9+ˑR�~��w# �ex��s}�|h� �8`��{O��Ƣ:�eh�)�q��*����u��Y�����"9ߍBe��f���m��q|�q>뺫��~���m��� rTǷD�ɔ���@Ei�uG��L��둮�f��1�qpB�x:0O�����������_��
f�3ߢ��d�N��P�����W&&Su�ݠ�z}Q���1�%�X��
���>��]��x����1Zb��{��)�c"�f�H��Ї[:���}��|5�y8F�¢h�F�֝?y�Qv���%�F�p�|\+�f8�g���V]��Gf{��ĨoVp��阢�Mqv������f�$ס_�Ӌ���%EFR)�vr��sY
�v���C�h'f4
!�R���-�|��
���df12u���o��m��|R%�����g������h�P��f������l�GpA����+�9��2�A-��kd��"�dn=���Ȕ��D߬��B��j �i��<o��z��U@~p��k�^�R/ƶ�����%2\�^	ʫ���~Q�`0��^Sv�"a���SA�E?��Bl���eb��ԑO�-n7_��9���	�j�z�/yj��Zw���s�O2��21l�H��d�������P��+Զ���2�*2�j#�jp1�����Xo�&4oX��H�ZQ`(�Ť(�GQ[����Rk���{L �=���1P˘�z��xJ���"+~��=x���kI�����!_�p�-02�=}�B^+j�3��IR���:����.���p�D���"6lS���P!59�æĕ�K�nW�ڏ�C��AXxj�բ���=�+���Pn�e�J�.�2rK���('7XfT�H�$<-@� +C��i����	xV6@4褱�Q(2H����:�\� yȳi�䣋(0S�q�NfQ�Y�uE+�x򝴥^���ʆ�� �S�J���%�YL̂�칦ax�Ӧ�%47~�j=�NVԶ
���c����%錂H�.��%_�����o�c����?-��݂�E"�U�����C4��������``�9�������/�����lWq<�YO�:˩�ߓ���]��BY�R��&�s h���F#2Ѯ^Z1����#ov��nI����u�P8-��'�y�4�G� �?��G)*�P�����d�֯��p��"��;� v����S$ }�,�vE���$Z2��Y�'�����kA	z����Bվe:8[M�SAv9��z��-v�;8�ρ������x�����+��j{�D�<dt���1���}<+x%�_����@c���ě�Iu�s�i��$_���A�֌��EU��ڂ���"�b�x���������9���b�s+ Z� H�<�Qyܟ[%�cyY�GB�H^AM�-�UW�+J	�yI@i�E����t���	 ��Jp�l j�Dԉ���Õ)��ʄS}�]6��"�?2��x��L��}Zh�$�~V�_T��|smN(�s� '�1�[7,2�|p�V��X�]e0��=.�����N��*����d�����6�LvQ�I���
X�r����K.j/zO��;.1��9q6̃`V���f[-�n#�zi6^��
EmA.v�m�,����q�)���v��$�  ����������q�u��Jsx�f<���)y�\�I�[b�� O�بs�^��F����B�u��H�h��-I^����VE��6�g�&v�5�R�ʉ�u+��t��������� ?li���1�9��U�gP��3�[���y����U`�"��;[�8:ޱ���(�z!�oW���.�P�	Lc0���&,����U0���{rg٢!+�[P�� }I.%�^�OD���ħ�ϻ�ܺt��W���H��N�b.��ƕ�q��or�����E��v?:���弓8�h�`7�����!�S���qh�oi6�QҢ*E���w�'��н���Z�ן,|����$�U��\׏��V��@��iAI� ����,^�{���,�*�RO��MR"��w7+��Ǭ��$L	7ݵ���fʡ(�w�K����b��~I������z����?�Y��0��(d�X`]�����^&\��Ը��ߖ��n��>�pb�����']�7k5%yf9�sʸK���%4X�Z��1��$�s/�D�M${<�M�[P�l��(�9 ���.AЫz��0%��V�|;���r���|+tW���U���ꡈ��̶g��#
�iy�Eާ��9@J޷��	qX�@�N�xXz��c���>�b��WӁ���L�{�#�j7K6O�
J��f9��*td��6�7]g�2~3�C����y�!N�%�⺤��g���[�)��<0��J���5�_���&B����^��c}�.�T7Bn*4�	�y�����?�`}ma����|���S���nL2r�sŒѵ5Rw�띧�K
l������������T�A}���K��3{��#��V,z(e�4��OՑ~<��JA��=b+@�
�ݫ�?T��x�B���UhR��> g)\z�W���.F]O��'J�Ζ~�<���a|c沭��j��sd�Lb��[���-/$U��YNy�|!��DP`�⁔�躇�X�rE�~",�X/���<-uU�x��#@��Lk��^��D����Ķ��w��t����Ҕw��'�E�[D=�J�k�5E�m�f�j��u=����^\IC	o�: P;G|���&�Ŋ��!��e[��
yO�Y*����Z�Q[l��;�>�*𣏕�{yt:��ysH4�m�8[�4\j�>�
��Ȳ��'�t~{E@qCpC��F
7/��07�E&k8�{t������W͜0�d����8�"�����6N�C�>��Q�E�փI(�1`����8h��$6�=������Q��"�
��88�h�H/FH�l9�`V�w爛����y^͢g��Lb���10��a��L��[�]�Y}����f3�h?�gu6R*Bl"fV���+��4�/�Ѓ)*=D��V�v�b��ᦢ����T.��F��I�3U��.k�Qv�8�c��d�s�L�2���aU\�K���&焦�ʗ.�޼&"=�m_G\7���R�ıE}F_�Nt�9s��M��sI�~�&?�p^:��cV���T�Z��.o���RA��A#>&W8�Ǉ�8j�{��,��C�(e\@><�;�� TZ�X���8��rt�L�G��8dO��w@�b��3��_��E��e/�$����n�]_H�>�&y>� 2���v�?�l`�j�]���m���/w0l��ˠ,��; �A1w�%�Ƕ���V%��G�b�TK��A�?ì{�S�f|4�=�9Ӯ�.ϏD�9�7*F�T�u��{���*�3�Vkm�2!���3k����ƌ��#7�o�\0z�s.��)�hp�������Gf�=���_m�X����{`P+��^W.g��Bv�"�u�����{�;k�t���l���37oS�B^�BxBв����Qx�����e�3�ᅦj�@sm��㱥��4L.#��G�k�������p��`�� 3�+�gV���8<�OQm�i�Y.������GD��7�3�t�΂�O�qI.<���׬�-��[��t �E��p�Z���q�b���At�����Q�����>(z���y��I H=�2��|<UT�4���
�q0���֋���n�hy�Nid�2��>$���9N����D��{i���-���}�B�V˜�3hgf	BC��jvvj��A�A��K+]�{�J�e%O�������ބ覌Ù<G�7q_�J����������0��E]Ӏ�?`�T��\ٛ�m�s���{7¤`	p� �������*�m�)���`���uP^h�^���=�e��ɯ)¤{�;��C����I�O�p�.A��,�O?Q��<12��	3��h�U��ZA�J���y�,��7e��:�b�Љ�������KS��Ȑ�uS�'���`�!'bn�b�x	�t��{��_!�77�+L>�C604��S�G���?���DFj�F<�u�{�z��l+�������t50��Fc)��>c��HcE���L��|��UF$� }�π������pT�f�O�{Gc�Q'�y�W����z��R����[ȏW��s�3�<��ƌ�����	Қ�[�I�� ]rF�R{��ޣL_o2~�2׻�5��>%���2P�^�1�q�hI����D`���uɑSdC�l#Λ�Y��6�������/��9Ͱ�*9�`���k�ܽ�+��Gx9���jZ�����y8�8���EU��Tm�ͼ�}���u��F���(�N�Q+{1���#��c?"����=�.�C�	f\����y��z�]�vZ�^�\a+�q�q��'s�d� \	�]����A�Ӷ�<����bV��������~�)M���k��R�lI�S{R*�&nEL��[ (s6|��}W3�'
B�[(z�/+F���O0���f����ţ���"�wA"Y��`L���d��j�/���)۽A�T�q��(�.�W�:���eRi|��$	��.<T-��v���®H��y��W�A��2S+N��M�B�"P��Eo����\9=�eSKC�0Ʊd?���C���I�'�+��) ��j��
eM
球��ջA;\uMF��, :���\�U�E{���^�m�Nn���g���o��jm�C�N�� /�+鍣im6��\��A?�T)���κ�ܼH�_ZS-Ƅ�Mc���03j�<�=�I-v�"��;tb��I�n5nf�)�Ӭ�dmu�3T����}Ԩ�;8�`�Ae����0��_������G�CÃ�K�'ìvY`�{���AV;��LЏW;J�|��Y�c��ҿd�Jb����m��X)��j������A�G�z%�p��Z�ŵ-J��W�b,`�����q�k� ��'8��|`s��B�����a�>Rm� � �#�+�Hm�j*x�P����N&ۣm��@�T7���xN�+�y7���m[�AM���p�]�zMxބ�i\��N��_PW=U��T�/\���plJ�"�����m�^S��E�kڭ�0`�)%Ѽ:�3ڥJ\+��H�"e.�Rv����wINŃ:_�E9�H���AG�>V���љ��jm>qy�����]Ɣ<)G�y�R��>dg�&�g�Te�O��5D.[�PJ!�F�Y.u&�f4����V��.8�ٮ{-��K�˙p����\��_�O75��ͪRs��%��f��x�}9� 체�ü��}ɤ6�N�?ff��]۽�%�ܮ�b:�J��ſ���Hl:���f:R����4'��P��&;PFoU#��n��5"���1z�t���z��zT�jo�4�u�a��I��R=7I��k�:-g�I�q�������D~��P�J�u��A�'�Ei�ح��ivًi@	�=��#ԱF^\���o�_�#���%P�&@������ޏ����,�效�$���c.��uiu�$��VF*Xq��g�i�X�-�B_�oK�u@ѧk�'(��N�6����e�E���H]��͉R���8j@e&x���$��u }btL�lm��T*��y�TZ�9�2��u�W �o+�#�#8h;F�$����'x� !����sQ?���u�^�}�1���s���m����l�"Fw�O��}�#��%�L�f %��!%�r$�Y��4��H��!Q�H>���-���0�ʖs�xltѿ�g�7���Rb�m�7Y�ʋ!}5\�!�P: *��@*�H�g�%�m24��Q'�U#���? 1I萹l���f~$�xO������K�ѻJ&��}WJ����F�3��v�Zlö:Q�s�gKL5�c���:@�%c�֮�2��	�?��[.C��m\�F�7k���u�L+覀Uauؒp��c�<p��& Z��	i�r��J#��g*xr�t�%�~4E��!./�>�7���e�^K)�oK�8ňFP����(�3�������Ѽv' �++N�K�T>�{�Fze�띗�XP{��&��#��q ��v�J�/��e˞��8c4$�K:W|����M2�U��FƄ��C:����ǽ��Z��=چ�v5%�Е�vo^
��c�͖E���,���]���@p1��k!�����i�q�14�B�D���t�~�;���eXgƩ2~�S����}R�f�l`���S�*y��X���sp&֮I��59L���_��H�i��E�}��?�f�}ae�ڲ�9��b�?	��Ͽ[���� ��\4�8��E�M�����+Q��'���)��}����{��:C8<�����_�;���]��KƂe��DEl^�l�qw"�l3�OH�|_^f��3�ԯ�zG�)�c��M�	*���q�"��*Q��4�$1�5���t>/SA+y�_~��e�MRj���.�������l;�@��>��@�/����𚣫m�|/��t�Z��PuuO��詻'F�XC��wB.�i+�P���L�����ؘ�u�;�8t�p��%W�)sO��ZwU�>���+^�ނ�.\�`1^�x�K%ր��e��U��x6�oK�G܎ʈ.��(]��W3w̦��,����u���l�\zͯ[�K��h!2�ڇ-@� y�M8ܨ������H��)l��������
o�5DA��nZ�!��/_b|'#w:!���>��D(MB8��'3��dJ�?dr��ІP;l�����6�,��8���f�_�����ZM)w�P�!���z]��]�r �w@|��fژ��`�'[2�����:3�_��{ :�&���'o��Լ�T~��X�\�wX֜1�ޚ�,�_L��X��1%�d1~��Ć�{��*Ho�h��v��۳MJ@EA�(�P�;����dREck�H�3Ba��jt�� �B:�@,���GQ���L`�Q:@�e������W׬���L�868��%C֗�Ḛ��-���	�t$��"��",�y�r�6�b�X��?S�>�s]W<G#�BAG�N���}Ww�x�ц4��$3��DY�A���ܴfvj�{d��(q\��ar~�ܺv1dK�D�sO$FߙcR�Swd�xíE2�r� �63$%�}�#�тI��[
���[\`$�_9��|��-N
|�. W�{� B�s�ؼoC浼����9נyMd"����=c;n�\K_y��t"yj�~���8�a�y�o��$�DD9��,h�C�9*ɥ�?ą5�lSᄕ�i%0�7"�{�
���H:���diQ�iX� ��I,m��E9���4~�J�A�6H���Cʹ��Yq�:J�-pKF%!�LP���>oa�ؾ��6�9I���y��F��{�b�8��POf�\�q�J(a
��sh�R�/��v;;$���;R�	^d�����|�n
:��c�moI��[�ƒ-��Dޫ+Ͻ�L��8�`~<�~�����:�O�˰�DB1���4<���lg���{��ݢ}�p�t|��&��ϕ�;7�6V
��d�{��-�q�Λ�T)�����JHqR��+ƫ�*�^�&ip����:�)�DfC_On���<���=l=�A���刕���0IO�H�MG��!m}��!-\�O` R���z4(��2]=/!���,���)��-��v�X�<�ƾ��^@�9b�dS'�^����M�����cBC,���aaJ��M����=��Q��cV�!�jemY�:��Y}o�G9r�YB����h��Z�s���kIũ�c�p2��M{����2���Hc�볚�
�9�K��7h�c'�^��v3��W�c�Ě�wƪRN�4���K:��x0���u$S/���c�7���M���Ѭ{!f�JĮ��h҂����*S��-�;A'&��o���>�b{��h
^�H��g㾧5�����'��B� ���㌤��۫d��t���^bv�Z��Д(��Mgٕߥ�iA�-��X	s�w�i8�P�:H���	a�'��h8?_ }N�h5�*��SP�87�r��E�ceV���tD�<�ڱ\O���p9#ȨQ8p/P��^��!ym ��9y��j�.�ҵ��5��Ѹ�����H���`�~Ρ�C��=�ۧ;�`�>���8p�ώz"�ӗ�'r4I��E"�	�uz��6u�򄊔�����Pf�#Xۃ�D�_�Ż�z��5�*m ��F���s������ PR
��+�!xԙ�v���� �q��ζ]�3�����ΰ�K�h��t�?�\��݅�ึ�g���%�=�R���]j�\�$�G�H�mb�H�(�+���/�
*�}�WY�'�/�ǆ�Đc�sL�à?��k.�\貃��`%�����@N'0����������ɑ�'2vW��	Xu�V�:�-��Juʹ�j��)f���A��_�b�6U��đ~B֢��a*��w�t�����؅�Y�x������gA�>�y^D9o��l�$��,�kS.�j��4�r��S.C��+@`�v�yUs����rְ���CL�ߔ�o�����l~� ���HCQ�
haA� +:����蘮�I��Mp ��%�,0cY��,,hA�K�{Z�R�Z�ML��s�X-\��N�㺻0	�Æ+�� �!���2s�y�:�ho����Z��!@�χ����K�屏�F�-!�����5�_U�<(�@M��Nm�X%U�����QI��T�J�Ǟ�4�v�4=����D��#f�y>��g���(9�(�Ւp �lؼ�t��sd0�W�~.!2���4̡��;� ��kU�g��䭝D`����O]��C��B1 N��x���/��#u:��x�zw���-tڙ����	]��"�n@��=V�F������9�橡�]Sw	d�OWԋM}xb�Ԓ�t��M�J�y^Y@�-�!W}�y�Q0��6V�A�|Ř�Zϳ�d��W��sg� a�H�r���9����N2����,��.5�ԺmL_�%�"ED�o�K�m�ZE?�f�@d���h�8�8я���%�{�ђ����]�Yw�j��[��āO/I,vN���B$da c5�d��YĻ2�\��b�]��G	�l՞�s��7�w弆��2�R��4�����w�gTk{�`S��3���'�:K0�B�8�w���?m���ڕ��Oe��xH+�tB�(�ө�Rf��=�]�)���!XC�����:tBx�
�ݨf)�i�ȧ�n�85Q�tk !<\�B��s"D�4�Л9&Òw#��=dO_J��b��t���ϡ��(��q����w[Υ�;�˫�F�-�����Z.E"�0�)F���-1�2<Q�tp���Ը:�@,
�gX���ݜkڭ���g.�N��#�_T>��������i"Ba����|瓭 ��ʶr|K�ހ���t�wd�XJ�^KíG�a������H'$���Mj�$A�R>^f�B����c3ct�����S���Yv6|ְ�r�f� 7���S��*�g5d�:���GX[;f��UD��L�?�L���W��(h���|�j��q�]�̝3'���y����o��X�g���O�V�B�����|��r�Їm�����M�ɃZ�_�Т)L?-ĵ*Skc����6�¢ڻ��v���p>�Gb��t��P���JNn���+��6�"Q2��6p���d��%/DIy���ضS�Ju�f�ַℕ��PI�y�)�g�# �֔ �-5Go�Xьd�)Gjh]����8�e��0�<�ue@���~L����#��@p��&�j;w�R���kN�"f�PH�V���N��?�x��$�E�9ߤ'�ڂ�ijo������$ʚ8�L��)'ŕ�5q�՟`_wDy����`*[����R|uǺ���'pe��VUJ>.ܘ)�K��du_(����i#n��"m�)�0 |&���?�2dBY02	W�~z�2>w�ՆX�	�q��31tN0ɑ�"}�~�G�ԸҾ���B)��`�k�!�cz������[ر�m���V󴻏hd/N}��ܠ%�a �Z�>]�����YoFdq��.�����8�}$w�\�~`?DH� �(��N�$������v4������Q��R 2�LQ���y�"���1u[,�K���"��^�yb�pC�'8�[�%�n[�^����q	��dJZ"�����+}�ʖ�\^��&����+��0����TzzB*�u�|a�/�H��J��#�QȬ���
�%d�?���׽��lBh!�j���X�N�h��Q�����#�Ȩ� Y�����\�?���|u����s�������U��A8�o͒i�RE8y$H�I��B/���A��۬��=/�� `��Ot�v}l�w�씕ȷ
,�Џ�0̊�MИ�q��cf�J�e~��*������͝"��f��9Еo�V(�"�)��N��G���d���u�k�_�+��,?�JU�K�����W��*b�$Yz��/	�����K8"�e,"m��Q�c���*T�I.��mФ���fWo�����M������B��<u��{���`Nk����u쀨^�j���7^6�)�Fs�nx�zp����kĆ+�?����� �e��� �p3���eQ�~ �G=����:�/�ͼg׊������|_��8�R�I5�$����hI�'s���_x�w�8����m!�d��R�lF}��Ɗ{�i��Gy�r�]�W���R�"�ͻC�i��=�gY|V������� �;b\�\�.B�C�7��a��c�B�5~�c������Ά���e�-πm|B9"�h��v',w�y��	rM.N�QJ\n���������j�VB��Y�=��X��<��n^Ӟ��-��5��]<�O��0�qS9o��9�U�g,�1
��kK��2�EM�k՞��#��:1��C�k�t��T�8�q�L���S@��J�y���uO�2�7��*�4�R_Y�*n*P�i�O2S���T܁`?s��e�3֐5^�_u��
|y�i�;/F��La�А7l���G��0��1k�����o�� d�݊i�E�u�����%��/��6�}���m���%� xx%}��
l��ZA5���3<@�V����8���E�2��f�k�%M)���X�t,[�W�bT~����9AVp���=����Ӏ���k�i��AfN�i܃���T�a�ӸLW���'H=f���y1wc��
����Ƞ\����@6/e����r�nfS����n��Y����Mק����Ywc	I.{De6r� [�v��/F�#X�z��v'�����OC/�6�ڧ����������aU>��NG`�/�ߵ�����1�D�g-	�>++��b	��f���h��4/#������pq=�E-��z �q��Z��NS-�/5�nr�
z}_�v;����4��� ��6���I�c����P� �Z��'	W��O$��#��Ƀ��0��m�P�o=�n�d;�w���Hh�V��w��G��}��F2?X!L5����y�&ʃ����bz���_�d��A��U�]Z�S�:_P�2X"Z�]iP�y�\@;�j��6]�V��i��e�5�cx�w���e؟;�����9��9��[��)��z�&����I��j���B�;��K/�+��F�duZ?(��<E� �)��a��e�+c-c��@�v �s���ո�+ppi�u�W}��1����8�8�x���=���Fg�V ��g{��>DP����o�7�牞!&N�p����V�l+�D&^O�V	f�k��x�{,�b�&�NX��n/�ә�<轃��!����B�4s����jcw"���Y��}����؄�w����I&��87�γކ�R���!����0\�ZtP�UK��	�;��
�;/���x�F�t;=�A;�w��f��s�7�BՊߥ�Y���,ZD�&�n]h9��-��L@����z$��*[ҕ��J7;A�&Ё��p�8�	�<�iG�~7ލޝKJ�o]̐檺�۰ [ӧ��&�r��Sc�'���,R����B'�&C�o��=i�� ����4.1�3E��?~$Kgh��9���p����n�~��ъ�k ���?A�VYg�
�;��V�K��.����O�����K�|s,�4���~���)'���A@���%��QC����.h,��5Y�^���J�BAg+�@	�Yo9���M�Υf?�v�=clp�E��/�����~�|���|����Z�^A�䆢��:}��ց�Ga�%"�ʢc��;�ьbjI�;������T��5t*��]7X�����aQh��-�HP�%�
�a/\��^���a4s�1�Uը�ʴ��`n�7Suـ�s�~�pǶA؜n{�c���s�=j-`*�,xo*`�>���Z͂6���Q�|����bv�ˎ�CA��D���54e�U�a�䠴���!
����F�!й�l.�������V<׭v��y���*�'�ƧPj~�n𭏺JQ����IS�C[V��g�Ƥ�+�8��.x%�[�\E��Z����`�q��q��赴���Ut��r��w���q`?{v)8�� �
M��_r���1%�&*��������PA`P��/'ot���K�PgDfQ�B#�ip:�d������+� Zh���^�H�`��[6R���.���.بF�^�&��Ϥ���~��8y�#I��a;y�O�V-q��o��@*�'���4��|	9�'�>���Kf�L.��ו���@�^y��V��G9x J���=#f'� ��p�\����n4`Cf#�H(�!�V�A��u�^��������<dS
H���u��U
�^�U�F��=8c�`�῍z���ؚM)��2����p��+-B��-S�+q)Goe���2�(΅#���c�H	r��l��%��E�S�~ڧ�n��y��H�ߪ8�"u���!#м�s�XiQt�(\���!0n�!'����̎�۔�rh�1��EZs�DIJ;-vZ��윜����"�4� �����;�9�j�UG�+E�?����s�NF�;�\+�og�>,��(@m�`V;��~B֙��a�t%������tu���y�6	8�����9��`/cE?��:v��_���]�="^�` �^J�Y��#��3=�i��%bz!g2n���;��������/��|�
����+���h�աާ0̌m��b�Q�m�oub�a+��;V;\�@W�l��|"e�Cfe�-�4� ��=_Ӯ�5���|���~I�? ���,�) ��5A��Z���0
BPY�]ck���:�J��G	�D�?�O�qݦ:O�J��T7��ny!"���3�&'�3�Zݘs9V�޽6��(.<?w�}��b>-UR4�!�ꞵQ��R�����%A�>DP�
:O��Y�7]U��*�@X\p��Cw�}c8^~�N��;e��9�@�"�_�q����N��v��-��R��X�g��wR�]�|J��~Ft�m�D��n��|�^�9��u��wX���h�έyc5�@6�"�B��p�1̉<�Χ�����i�����o]��⯸��W,�l��鏮H���&Y��9q3ߺ�r==�?�zNl�)�2��iƋ�Lt�2ȶx%,!���Ww�0hH|{�uz/����)�J�AL�@���h���~"��Fz��;�!�3�o���^�=���IF��ʗ����Z=j��S~�m��s��{��������J�� �U��T/anѳ��/�sn~���oi�VZ���:6W�uAURMy�4�B�� ���U�j������Ɖ���>\e��2>�l��W��[�Q��9fc2�r�`�?���R���qrѰr�Ba��b.|�Ԯʨ�)N�jwiۂ��d�F��e�[N��IxE��r��}=^�� �7:1`��٥i�)��hў��v9����D�n�a�D���z�8Ɏ�0�/|�j�(�βR�<l�N�����>8���tK�nnФ�1�6�
-
�����7�C
�1�kV������pf�7�@��DPM�ɈK��;��}��5���ٶ�z��K�b^"�I���M5rq�k� �	Ao�!�����B�Qk#d�aCRSH��!�P�*C�(� Djes˕�K� ��&kIM�J	N�c��SLB�T��� �m��#���T��[}�Y4/�A���,'?�3	�	2x1v{ae��}��Y�a��?�y� �,��O����'U��6𺘽�]8�H�"�w`1��(ej�'�l�ċ8\WC�lS�n�ݶ<\�龝#���Y:�	OmPSd����M���1�N��g�:��^f-}O_���G�Yx-�o�ё���ǋ�ߠ�Z�Ϛ��:�T��B�1�����M���4�C\��͖���a#n"�7���{	0	{�������ԛ�wK��l�+:��3.�۲̋��ܥY�������s=%u�|��0]`���~�@��� �[گ*�<����G��k��r�'	圫�ܨ���P��[g��y�L��Sx����زM��8ݹ�0�� �Ԯ���?&���v�D<�d�/aK��qN����?�<�-��6���0��a
>�A�:N��$
����%�D�8�7 ���sv+�Hоv����a�j� ��5�9����U{�S6r�BM �(C��@��mZ_�tp�E�Z���2\rK	�q��X�m�$��7j�w,
-�s:1�0좥�V�}a�T������%K�"����)�)_��	�����tD��i3�T���pp�'��
������7�۱l�%Щ��oH�� ��<����&��_��N��X��T��{5�z��A�0�޼�--Hg��%]i�Q#W� _~4�[���X����L��ۉ�Bb7 ZJ�M��U_�����HR���w����g㏑�^t��e���j���Pou]��ī�ZGet����sPd)ŘZi�b���ӎ�Z!M9�c�����I�Zt�OS?>���b�t���&p��c�H�����ڿ�]�q'�����h�&�yB[H���B���@:��W�|�%�>���/�C�|�F���a`ǯ�/�R���{W���	�$��o>���Mp�CO��b��o(��K$̝�	"�e�6o�\�˓(�٬��s���a�FQ��iT�R�Z� ���{��6�� �<y�Mf�%�ηm�T�����h�dMS�L�[�V;B{��Β��`���R�q��,��8k����Sc��Z~Q�����}� ��@=�`�tChl	+�wM����!��C��m1j��fY��Z��@��8.��e�x���tO�g�X�^eWԺLmI��RwK�oP>{����jx�X����Èq�7�-2�𰳛YF�l��X9���sI�T!R�(���S��?�l@F�y��N�j����EӼ�o}3-���J6Zt��|J�c���'>�8��"�ߛ�)��U�F+�{��S�Vz�<{S����~�
�����Q���`>nZ�K��ݐ�O�"����1�=�h��X�a��_�(��n%j��8����XI��uίHԑ/B���k�5��7��|��3Q��g��	T-M'q'
#����s� �~yG��,���W��$���y9>��e҂��8f?JX���u[�u�Q�L�wq�G�����x-���И,Q��<s��ҫz��6	$�"��K��4�K�NlM�,��x+�l�}��A�s��9J{�+��|m����q��v�$��P�!��C�b?9�wu��������j2��+#	l,~S���S�'�'��d@�܀�^uxU(��vN5�c��`�lP�/�A��NŇC�b?�����J�`Y����Ū]
,s��:ӫ��ԏ�l�V�=�н�ss�C�E[� �^֨���0���_;�~�`�a�,8M�]����!񲙌��>��co��t��>�2�ªR��,f�Ǔ�0�\��8��ٽ3���{r�T���&��'����K߭�#�	0x��µ�ȩ�au���W�p��n�P\��1
������.�t?������.o�O��S�^�'||��9DG�L�� u�]�+��0�AD����7�Jjz5ևٺg�ڨ����6�GD�r��\�PXz}b��de�^��ך�XOywm	�\��2��dL�-C�zg&}b�w�5d���$ʯȌ��!�s���*�o0Y3���pg�9��f����P����U�E����O9�+��`����=:����<����`9�; �h!�7~aָee�+��9�CD��S�Ϣr������)��9+<�{\�%ˑ�� +� v5�V�.��Ѽ���V��^��5&�����5��j� Q�����;�9�V��A��)�&�Lv�J!54{�=Ҏ*�(X�8!�:�NsBc9���WsĊ�$H�C��j�s��+�{��@!g�w�B���f��>B2�F�Aʿ��1c�6 hDO��+�\���n0��Xq�8�Q�ν�h��2gX:N���\��ʡ}8�O�	��C��tG@�ҷ�bn��7����{��� �+��k	�|�_�V')�{lDhG`O�FI��%2��l̴���#��HS��'�|����B���es������2_� ��/��OQ�zZr����_�)�><n=���o䵏����MS X�NRJ_��2�	k�Td��p��nt��K)�����r��+M��v�_-D�	�Z����v*p�T�5!r#�$�y*�Upf�Zh�/��qCF5^a��C
Z��	ySH�В���L����*4�@��?ӿ󉎔�8��4������Ƶ*2)�h����<����8L��m�6H�se�[lvY+���IC]2,y0m��?KlC��xa�Wl0�řs�L��t��/ݙD��D�K��w��=6����X�-��G&����}�K+�q}����]�P~�ڵ�?p��R�����ŷv9f�2wa���QN��c������L.?@��n���&���-��ޒ�R��`�m���qD0yA���a�`��X�`��r14`���#��&������̀�t�G��"J�����gL��
t���b&a�,K��Pd���oJ�U�ŝ��2u�~�ZaA�]��I����_6EK?ޅeA������Bͫ��%k��w�xP�	����&Q2̥��DP�c�N�#rͻ�bK�n�
Ŕ��_���n;腅�����SN
�ٷ�v�[( V� u�'�Lqh�J�FB��3`o�03X��_��H���j?Q~�j�Ze_罥NX�����"�h�]ox��ґ]��z�,���Չ�6���
�~�)ŋI\�җ'���+5,?M���-<���F�ti�A/H)�v��#�؉y�~���6(�έ�e%����(��Ddb��Ym6Tz��%���McmTV��{���$��V�7��o9��:���J3����6�Z����$A�D~�Sc�"+�U^������
S���w���!R�9�1��� [�<�d��������S ee6��O.ž���c�=�^��l�cjg	{�ՙ,CpeB�3�x���O�y6x���An�ͬ�U��"�����(E�̖��
�O���Z��_�
j;��_6��X��o�_ d�;�ܾ��:�B5���B����������zv|0�Y�̂��]��� ��甁gr�=�hI�k�`��`��a���!�Q���R�:E�K��m;��Ş,�=Ax��V���pS��FeRQ"rc�!s��	�^��ʴ9�4 �g�MO�3E���1���
z�r�p$7d����$ocؒ�
��p�)E�|l�r��`�ݭI�����]���a�M����Ѹ�򅺩��%��d�r���y����ƚ�l+���M�l���c�4�kcF��"#�%�-;�('1�K�rL��9D���%�2S����i��읷؞��y.�>%�e-�؅��R�$M�C�.��gZִ)!kzz5YM�rM�)*��c�F>�'k,��J����Ԗ��#�((���dV��۾g�BϚ���!@6ђ����3�ۆ/s~Hv�"�΀�������Dv�F@(Z�2��q<�'bf��Ub]O`z ���v��`�`W���G$��-��Z�4��2L��v6`@ �Д�c���� �Z���HN��X�'�'t�	)�vo�G�(W�3��G}�{�,&f��FJ����d�j]��O'%�Tv쩏ySP�.<֊j\	v�����(��f�In���|.j������7d9rϸA(a;�n��w����̹y'��F,ۼ~��������-j�"Ap��-�U�V#�Er�0�dK:�Ö�*q�u��|��ǳ��X��%�f����i�v���Sİ�d�J��P<��vZ�E0Q��C���:w%`U�u�)Ą���c�m �c#R ��/<o�Aj�`!k�ɨ-LU۱���x��!7!u�D}�C��L��U߅mw�l���N��N���d@3�ȹk����D}���e�A�g���84�p �o�k��}�\�����hE����yE��=v@��)Db$KyZ���BN��u������LzAfa_g�֖Z��+¿���M��uN?�T|,f����2��4Mt'��?�=��r�l�T���V����֨��!���_y�\�w��pf��[��+���~S��U,WF�w4sxs�l	][�4��D���ɇ�TNȺ9\S�E鮱-4(��H�@W�>N�T��Ua9x>�~�7�Utc$�᐀m�U�#Xރ^!�c�躥���8z����
SQ67�@� 8{E`A�OIwߠ���xZ���~*߬癭+=���iV|�"_��%L9|�5
�`�j��>kw�E�����s�����g���ٰҸ�A��}[Nݐ��#Ƃ��<�Z���c=�"Kv�h{�����Q�xp�Z���8�!�Z��/w���A�Au�2��
BP�[>��<��CXT�)O��H��������b0h�b�<�\m�栆���5�h��N�q8�[�nr���f���YG��R�X�������5Q̹2���eQb[�Hva�L�t�`�^,���H&[ PtC�K�i��_���&<=��N�0�ik��W�g��k�{@м��R�֎:�v�[z�b��:V`���/�A�L��tQIM�
$����z��#&��D=i�%1�~!����&v9�D	?!	�;�c�'�2�*~L�:�@ e�lM�Z�$�@u�;l^���=81��Kb��u�{�wᇀ��!.j��̃�a��jVq�Z:{|�f{�T,u)�p���LX��&��v�`�10��K������LJ��0�°J�k|����A��G�t�p<����^���%p�q#(�]i@��t����^�*��$�+�M���	û>f+$���H���_9擝�b0�RF��.wi�i\����/�	Q����cZt+6����0#�n���~1.x佁��0W�5'�d���~��#�zf���΅=�$����Т�rH&e�O�����A�*�<*����*�������fpc��#��q/�W"��=��׎L%K1���լ�g����0�/�]B[����N���Q�����d��N�.�PP+�̅�l�>ݵB3������7��a��{�Ȑnw���:��?�z���OS9P�{�#?\ĈP\��;��`2��?�Ĭ�p�����y!|w����[aR�x�)����REˎS��,���}F	����,�{���i���U���nB�\�U8W��w�9�1ѵ<������y�`o;�����0C|�c��?&4����S��MM~[�������ftm��j}�I;��g�5��I-�S������P~�4ɜ�	:�K��K7`�$vQ���AH;;u�U夳�G+�9���m�y��������f<�׏mb���3�`�̠F�c6�.�h�O��W��D�fX�6�d���h�����e�O�"�kg}��и��� �J2�q����~�>|�[1m��]���"F�s�P�X�P{٨���T��z���e����JM������@�R4���\��Zh�N}Hn�(J�7��1�!�^4>J�qd�8㥢;�b|��6�8�4prg;�N����s������r?/fl�Df�x�e�!�8��>Pvr�Rm������m����7N�O���O���M+ק����Z��$E��@E0+#yg�H0#��X�Z���J��.�bIh���Dgߢ(S_��9l��S\gK�}WҤ2��0Yޅ#����Bkb�G��FS�p*ע,_>��{� �43-�в��r*M��\r^���7�H�Jvq�Ad���<˟���N޲v�`�G /"g���ڊ���������I��0�� �:��h'�f2��E�cm�e-�*<�����<��U���m����v8c
 r�`<�rV��Q'�DފhbY�\8��ǲ;�����Y�TFK]�Z����͑����gW�~JY����E�H
����������Fa���S2"x�H�{DK����
d�D���i7�����`q��	?�/��)Oy8�٠HʺU���aw���P;��H�LvS5t��Rv����e�U�G�4�x@���U�>�aC[7�ȗr�o8�컞{@ʻ�h%���Ӻ�y�G�����u_=:>��#ջ��N��0'��t��0�S�^]��4S\5��m�[��)e	��������!"
��7ܒ�l�p����[�ʹ0��ђ�O�G�-G{ s��Z�i�:c���p�f��A�TX�e+��;�p�`�2 ��>�WL�7!=�Z���Ot�-i��Đ�j��x�=rS@��;� �+#�o�UL����PW-#o�{�S5�E��kc��M�Å�s_vj]�8���B8�2��"�m"c�%�5����ʇTRpOu����{Gq��B�!�q��)� Ԕ	���/�k�{qzj��r	3���$.���Q�b��My����q�]�����%YL+���P�љ�����`�W�!DҰ5�)�:��o�?��A
XEPf�>G�įPҜ6���2��j��7�"f"�Г!�k��\R�1)��b�U8fѓx�{����()'v6E���/��{m�Aզ��؞-/��h%�
��{^[3�w�������~ǀ)H�͡���K3�h>}��1&
�8 4�|�+�&Ϋ���.mh��Ǻ�8_�ĽjI���0R���*S�=�O^���,1���C�'�Z&�K�G�:�-��3yǴ�I�'���==d6���N?Q ��Q���a�4j���6�b�R�k� 0(>/��sJ�u�6��2��o&����D��LN]�2�,D �S}�����o4�K
�U���t�M�K7��N��2�9��Q�;��7���V>���	�4���<��8���[��4��������p�����<�	��B�����)�d��fQEkʽ��e�� ӭ��Tg)���G^���A�O���Z��F0[�7m���l��/�%��Y$�%,V�4��BA�Bg�@���X1d�+2�C�~oh��]D$�2a<}��hZ$Cڒ��<l���^�^Q����C��� �)��-�I�����Hn,Ⓣ -���F�p74:5����Aa�������˞� �?��ˮ�kr�<t��w36�S��#�Oᅼ&�#ȟ ��5�4
���F��>�4?�����)��]l�*�I�7���(1���@;r-ϔ�Z�����𧃸�S����~1����j���xx�&ч�l���I����R��`��Vfv�t1�8Z\��JO���;��_���o����{��pi�-]��"N���~�S>�:�y��1MĤ�Lr�j�� �4����V��.f�|�s�.�\a��&�r�l4��@	˯���^��*�	u�1G�	� ����X!�a3�(ʵA�Ul#hC�|���8}��2�ہ�- ,�N\�H�*eW!� ���9�<���8��c����XK7�S	��i�G/be�e#�����q��{]U�xr���,�6��ӐM�]gщT'/uL�+�|V���=e��@���F�0�#c�ϛ;Sq�X3�߼2^�M���K������y�Y�ŀ�U��)ED.�:H�2$ߎ�D�V�	�z�s�G2���ʏ;k����߂~
�q��s]TK���1<0As�H�8�݈&�g�kT�8�y=g�y��wek+}K�2(�>>r�@r��u�65LKl��T���w�~�YW����7����g@��Y�m�?t@���o乮7�)5��W�a���
?cLo%����aίV��0���@WS���v���_��p�n�!�a1iB�� �w�����5��VU�wU�����{���E��W�C�IO�WR/�=u���Ӱ���ӵ���U�1�L��М�Z��N���޾��� �ys�$n/�fHAq�d{��+f.�{��2$�	��h!��e��W�kp�)��嬼-u��N�7��\|~��z��#LHpt{E�����h���{['�,Z0��Y��������_�X|��/�hIh�]���v7�<���xB�
/�?z�nɆ#8�55������1�O���"8��˖��)!��pZpO�O~F%%0<2��_N)ד�.��Zͧ�Q��25:��gK:p|�v�Z[Cc2"���{hz��ւv�����g�N��6Ǫ��0���)�����g��AC~|��S�]?�(�<�2|XGf�gf��b�]�&]��p0��h�����+i���������S�_��}�٢qMQ��|�r�Z�Ov��@�3[�k�0����D.*�`	ʳ�|��LM�W'������|�Q�V��[r	�
�1�0��f�2�xn^(w%�zl�Q�]r�V��1N�R��]�E�>����'w��O���s`��{ {pP��p�[��n-_�t��l�������[�q��H��	LN:��ށ�
���H8��sI�5�5:X�@!CW7?��\4�˙V`�jBA`�-�������%�����gy�ż2��G���'�b��.��S��=L)�r�G�U�|O����_�`b}r2�xPA��j�W�XX���`/�r��۲���<��|������	��CH1�+tT��L$���F�.�~����H	����$oJ:�q��E�����9��ѨK��[*��db4�lfo�#�f@x�����!"�'p6 ���9�R��Q��W��K��������U���ٱ�\�-k]��>l}�Ap��#���!����7E��'��g�F�Yz��݈�w�)���~��(�0+_>�O��΃������JN�nU��O1~��ܿ��:,���U�q��v���"�݀k���0�
��}UD�}�i�[�u]�����l�-u]o�2+�����\���&
&�n����`��r�/f#��]q�BNq�Ly�2W,�r�c'����[�cP����]��{��zGԻ��[��ڢ�E/��y�<V��/������#x�l-$/&�Q B�/�2�4�S�k������̄U�V��C\�4��΢�����㋶,�X��ik���R��'f��+jf�rP�}��*��k<P�*��҅����q��o*�3�}G�d��Q�9�M j�Զ��4��9���Ћd� �8�S���$s,�Zx�}%&��/Xj)iņ#Y�����7$?&	"g�4�a{m���l ��>QN8~M����w�|�vn�L��u�ά��[��f�`q]�@Y�rf��#X��&?���5��oh�J�6˷�z ��Q���Ȯ�~tο#;�|���ԿSXqs+j"��f�9j
ӬIm;���&֬4 �V#�U�d�ә�(p7l�|�b����_�g��Ss�G�D4�
d�9U�}~q>7�����s�Q<��܄vQ�M��E���d�q��`/Ud�E�A��\�i%��
��R7�q�<݋����;փ7�zF]O�C[�7�8E�*;Z�'��t'�3z�z�ᓎ{C֋[�8�۱�(��b��%�(�yz��d���n��O �/8�9^��rUU�ؗ�Y��T̳��œŨ�$��0���N|x�,��Sf��8�a���$bzD
�&� 8���/o�v͂f|:�E�MeT��ᢑpp�Ϸ.g��*�����Â�\� ���%)*�ο���٬��8/�|��[���=d|�^n(z�N�(娭0X����D�{#H�<�:����m� �/�e�enV��Wh~�d��p��G�<��7��U."���h5��B��%ދ�zy�|���V�č?�g?[�@~��w��Ƞ�6NEf���;�ZZF��%��'��dU�����#/?�[�KQ�j�T��t���q`he:$���1Gʤ�T5׃:�V�(����#���1�]u���P�J+ag)��ʬfr������:}�G'��$�ʯ��<ڞx��ݎ�����QE1M)�ہ.]|ހӷ�;M�����)��:��ED�S�Q?��A��}nzz�st��Rdz�x����Ӝ'��\�y�ny"q%D|5���p����}@߶2��~�f�����w'�2�S���f�l!����C�mL�^�EZ��^���f����D��NU��1W鶒՟�I"�SȾ�;B�!�=�
+ ހ^Y 0��	9W�%��5��*�@�6~jYQ!{��΀.�yF�V�'�;�WE�x#,��	k�v��f�ܑZn��4��y(U�\�Km3�#Ȑ�{�?y�78�l׎*1�82��5�;h��j�M����>����#��\��g��XWN#��ߺs����ߑ2���=���}���2�	�F��Y��v���Uy\j�"�y�uvh^v�E�E�͋i��v�=���j5��ԸU��7=/��6WB$Y�24ƂKDf�	�VV���,5�z��+�����j����3{���a�ٖ����!�BGƅ=,qY�lg��O/ ��*EM���A���,hX��ȹ��^v%������A��/�s9b�
��+T�����E��g�3�U�3�c�3C��-�N4�N�rˌ�E�0T�ۋK�����bjFl���gU*���v��։<������(�Đ�.�����/�<�7<��f�BO���a�a����I����x�;�\C�6����N���3��n�U���I�����X�LV�$J��,��#d�ۖ��q�s�����_Q��k�φ#���Aj'W�Y�Z�Die��-��dc|Tq��(X|,WV���+h[.�,_�݁Imc�!��P	���h�_���[}�� ���cR��Wƅ�^�}ӛ�|�x�m*� >�����s�'��1�<�>�R���$w����#�v#@�h��Jt��%%UM�:gC�������v�o�B�@,���yaTu`ؽ���w|#T�d%���<�R�_4߷�u��Ku�ܿ ��sQ��^};vgqb��BHYp�e���4�$����f� K�ccbZ���8a攺V�\Ca�Ձ�v��W�?X�7(�u�o�$\L��yd5C�\��@��{t�������j�$���/� �/���B�������Q⌔y$�_1Z+)��ǘ�驕��w���OS����@�'�פ���ʮJ1j^0{�?�>��Wh·�z?�g6�����;0�;Y�?����8�z����:��B<�_������+=T�.�J��je���f��bbN����Hs��������e�OP>OԀ��U3����:�Jf�1��>�C��w*�.�[�ʢ�fC����/ �ߕ�H��	0�N��7�es|p�MNmO1*!���i:Em��ʫ(7�~�F�,�&��1O�������3N���ĸ��D��_6I��͛�b��J�|��Ӡ	>���4�I�z�։�x��ts^�l��φ��C�wÒ<F¦��A��?L�~:��3N�Y�� Uȹ�~�����F/��)D���'���T����K戀�\^�����	W�o�����c02Ll �H왹Iz���"��!ӄ�l�����)Z!vz�2�V�L�p�%�����6^8���|FhjB#�(�_�&� �X{��@��x=�-%@����>��^d��_&�>��5M,��w
��T��.��@I�B�0ª '���J�J��`<'ݚ�];Yǁ�n�s�p�a��: ͪ�sb�����VU|M��|uf���+���>�Zh�?y��B
h\�����z�i�a� �-�
��Yi��Gf��
u"�R\�,=��weZA?[�%�<��r�
�I�HH���y/��]ǟU� ���M��g�U6'�n�0 `��:�W (����R$�X� ���\<�N�+4h�U�?��]���'�Fm�1�;��]U7N5�^���.J���aW��S��]�y�vv�����YO�F������S���|,AAi.��g]2�{z�u���,����Ua��u�'g��#����'��&�xbM���;�t?q͢�ԺZ��Q�h�Ejו�Ŋ���	��L�6�a������Iz���.�֑g[]���)d��D��G1y��d'[Bݭ0~4��!NKT�W3�9�e�0�R 1h�P��^��2���6*�����z���5tLu�B���I��d�6d�T�!\�\!Z�������bҨ*��I���>pz�u��!��2H���b�H�6<`׃+*j��� IM-���t,ٻ��\���U@j:���Td9�P~m*^W���,�Z�2G�7�s�A{;$�T�r#��m�����|ً���'\�VT�,�~�5�k�6-T3��uᝊJ���L%�7H�U����g��(k�CӞ;�U��UN��o�S.b�*~mEϓ���u��8Ή��,l)�5��'7��&'Tƒ.�^���&u�*
����œ�S�ΎY�c������a��9',߬�6e�v��rXF�ai���KC�a�W�	��)Yv�,��ؼ?�ྶUe?�hYㅠ��!r�f�l��h�yVZ)=�PV�c��Ͱ�Y�1��&�A=��:�7�*o�`���cKnV1��<V��M���6�l����z��e&2��/�a�k���1oދ���cTz_�1-�B�����}e���R�RBsA9+����c� ����ؾWǆ��v@Rۇ�g�L���@�����̦L��z�M�0�E���v,�
���d`)G�!IJ��"��hGSh�w��9���Xy�m#hr��kl�B �.�A�,Õ��e_$4Xrz���,եJ����:gA{�:��g�1&V2^v'�޿������̎��=s�Q������(3!�r`�1@m>/Y�/�G�&��M�n��W�]uծB0G�G�?U��_���S%�+a�"���Ox8SA���C�ޱz!�8*·M�c�����k̄4��w��[�>WH�ۇ�6�D��-��Ld�����M��"�u"�%)	g;�I���d��*��8=>�O�@|��-�T��7��,�Qq��Q�=����R�� ����D�!�;�]��%��ʜ����-�W�oo@�8a$�=��õ�����~�}�ty	�q�MĮ*QE$%*3"��Et�a�<}�B ]S9�:)�*M�jK�9a�Y1�n�K�:e*��̩v���k��ط�8�x>RD��6�$+�Ð�����C3�-#ݭ���K��)[��m]�Ƭ�/ds��Ì���l�ӘV �E)���o��y=7eQw�P�t�^�rR]�$�kʀՁ�@��GŁ��T-�T��Jw�x�E�T|�#-�� mE1�w!��V�o!,���<g+C��h����IE�]�_���TP��O	`+���wK���,�` �n2\����*���~Aef�w�!) ��N��>�+��;4�!R�b��I޴��ڤ��������.��[��o����u���-n��> >	$��P�&9�dF}��I�0I.�a^�*���f�q��ޛS���AJ��#�h�U)f#�)0Yݓ�Z&O`�i�^�;���n'�lR��@�	������H�.�E���X.)&{GoQ�J9�����,_��X����?G����:F�`BEam��8�9#�Hk���%ɪ��1it����]򷦦����p;�����Ym�(O]>�6�Yp(|%x]�$\�d�L&�5�`��`���&g1zҷ�����H�eJս46��0|����z�)�CN���tc���(@���ǋ
s�y\NRvP"ݐ�|�f��gz�_𚢖�X��ۚ�*&2�-]h��=r��gSm_��)�y�I6ʆc��O��۵��g��bP3�x
I;�ʡ���K� ��	:�a2r	��cx�3ά� ���r7Z�{e՜O�s_�
��eЋ�$�!ob���1q�v�]q�W㮈�_���퐅�S�gxΒ��m�ی���Y��#���4.�F`������Qo�ep��bZj��}r��hӤ 	�Ib�'�'B�]J)ۑ�H���]a֟��b[�`ō2����HP�=U��.gy�qtO�(��6 ��0�}��
�5�D�j�d�>�a�����*=I���Y�,o���MV8�S|Wp�C�Uc��x{7bg�LQd\j��	K�y+�Lt�T�y������FG�s,�k��T�VMH�g�:����Kc�!46&d�%%=p�[{���%�s���}e�1Z��G��ɍ?𡚆(q����ɢYb	#:���k���m	>a��,�P��n��$���|��)X�>#��.���k��3ډ@*��G�"�d�z��t�ϳ@[y�=}v
�$��ݢ�
�������J��N�Q�{p�GO>2��'�)�V��̆�P�\��:�E���B��U����b��k�&�[��IP�`}qU� UP'�h�<~y�2"y�ꈑ&s77ټ4W�yL�![_B�:}N��Fq�0� �<7JD�y_����g�,�HXw��k�P�`!��zD�yE"���P���vX�@g�0�q�\���[$^3��]��V|
=C�
L����=ܻ��G{�i=
�l~�|�Mŧ�nw=Z��s�Ԑ���R�*���|kJli��E_e�(ۣ+R5�3�=>˃fӱ��1��A�I��lC�o��p܍;G%�ZKub���	�?�蒣oW~�u��݊�kP�1H7�q�-N�t�����Q�
�>L&�4g�XY!�d#��]�a�O�a�ؕZ]��
���B�p�Φ���SK��Wܖ�f�_��]�ͪ3�.�kR��׀J����h��ǆ��AI��qp���0�P[Ht�(3�	�zDv6�4菤���ݢ㧪��9pf��U�#�`�`�paSL-۸K�8v��DJ��j2m�*��%)k��������aQ��fX�X��@��"������F�k��k�5Y��'jz|�WYq��-z�3qB�3�l`W�w��=
��ʎ/	=�-)0	�C1��U7�"M�w�f�*څ���%O����/�-�yޠs�}��F��LZ�m�P�,�	���#󄴡7 4As�#t��-���`��z>�L0hf���&E�]�����g�u��_n9j��i y�w�Q#�� �ź��1�ד	68�`]���L[��Vǧ����@ͳ�[l|�8*�{��wP���x�+�EL�J��T�K'uT��7��Ģ�����D%n��P�:���o��Uhԏ!�H�r@��H�uf2E�<r�0K@���bEM�i�E.n1��y���cx-W%���Be�"z5rǓ��mQ_{��\���� h��+bV�7G����G��eM���"�����g#QI�X+�G{Τ[>r�ƺ.�^\�e@��Ց?��M �W����3���~#cqpd)��j�`1R�/�؂��� �p������o�$J�/��\ 3Zh��k�zlx|�[���|W1����..&MH���+Z�%÷�Ӣ��3����)��ua�CP���)`��s���WT�.@IH�%3Ɔ�>M���8(�o�<d�4�!'7
�oa��@VqC~[�����SR�z��)�7�9�� wK��[ӟ�\<�9� YF�vj�l���E��@j�O�D;�����'��,s5�aDFo�4�[�SU0V|���<�=� �5�,#�� :ɽ7v$�}�*���}^:�cO�ABf�C�Ƞ�N���`J~{\�bK���i�Z�K�>���5�����Ny����F?�>�la��nH��O� �r�?"y}���V�͛�'�a����ꭈ�&P�I^��ک-x�­d�W�����r
�`N��!�C���xT���-c�m����\�u�Fa�X�&��-����;yt��?�l��7����i"Aؗ]��Du_@~4�9g�P��|�",�҄Q�6��7�x��a��F��'x:�
�p��b��V��-�5zV4�}���)[��9��9ڡ���� �q&!4wZ�D]�0�m&1�@��I�iu��P��x�C���g��_]9_4[���z�����#�"*��nB;;{�<�6�����q�p[��8�����:.*���a��Sa[OE�߾�,ӛX��)����@�ƨ�;�R�}�j�4�%�)
ִ�t���^��֯�&�{�"JL��d�|I��"m����K�g1���ꊸ�$i(�ҵ�s�4@��TC�]�2a�b�#Q�+���>̾�di�ɆF��hd.�h>��@��9�:���q6xaw� �+h���ߦ��V��jH�����`HԾ�-A�2Zq����"x�3�;�|Nl�&fGne:Uǁu�f��l�p[#u۫D`�g�/]�	�����t���5֪uS녕�%&���gt�b��d�`->�6^�Gp�r��̇~��z�0��6ȳ�8=M9;L�7�\�<��{��[�>`�G�1Y�x��3y����E�� Syo�pv!��a���5!dU�M�8%�E�ș  !֓
+���4����{�n%�2���%���"Ű����g6b��G�;���%��c���^�/4D�-Z�LPy�J�C�{t��7���`��ڍ����n@�A�hlB!9M�M:%����i����F�!HFm�\B��F7f?�)�q���K��tԨW��D�ES�$�s.��o3� z����` ���p���$������D�*��U7�G���KM��W�V���^<��Q$L�O�~xZ�C�@$ ?�6��{E`��4<�JR�.�qo*���$m�	�;R	'�V�T rh� ��i2|2`�Ng����Yy	�>z@�oT�/�N�|a3W�;:"J&$�N 3�*�7}i���8| �<i ߲���KGx'\~���&�}g��=`�K����4�
]3���-u�Û�.�4�G�i�̂"5�z;h��F5�]����"�f�EƑIޚp�{;9�٬�k�Cj<�?Z�a0;;a��ʗ���*@�7���"֭�l�L���hCy�G^s��i�.V/�$,(�R�h<W� ��[~�sJڧ ����@
��i�nh���V� _�Sz��7n+�&Z���x��i��$�;p)�q��hȕU�G�4��� B�������g�� �_)F5���IXX��,��Q�š�~��ʲ���{a6)dq�&G�?!~�U⥋�Լ�,��x�:c'��Y���'��s�yR9��2�ƥl��4Ҍ�TV��=�.�G�}}O��YD�a��\y|�k�D�����4�)B�j��V&my���ܙ��3p���)C�G,ߓ�x���U��t-�t�Rrd��O�6��6oj�G�8~�̀��?7��e<�����=o�1mu*��p�C;���x���c��eGjVd�舎/�,��ڑ[H{���-�Ep�f�������	�ZW�&���s��:I�Ag��X+B�cO_~�]�}P�Xl���L��e�.3����T��ό9V�W2�ǃB�֙�b+Gэ�]�)�gV�	��T�;�.бPk�Q}ڟf	xY���'dzL�D��V&��_f����m\��U}�BK�z�I��֦�"��(H��)���a�$�U��W�&`�ȹ�j�[�<҈<p9�F�a�J9aח~'3\�Z75��S�6J[�����e�W~��@���n��W�h臈���"�HDȮ�,v�`�*tL�5��Uh��J%�C^�+J�h(�.�$u��5h:e*U���J�}�2cO��Ɏ���l�/��������S��f��U�O����Hp�7�rx�T��\�2$�R�y�D"I�Z$�їug�"�,��뼼IѽeH�"���=MI����Ԯ����$a,������tm՞uaՙ6��X{�$3�T�`�2W����oڣ@��C����e��Y���Sn<������V��&S��+�٩�"P"��!�t�r����U����X����[�5Dih�9��c~���H�a���ܘ��"�u/L!9z�	�S��_�dv�ջ�z��H�x��ӆm�\s�ȴ�廆P�S8K�7�s��Ş���O�%,���Ka���VT��54��U����h�(1�)���e��� 
1�=h�ScN')���[żMj�����3wx��0.��;=�f+�$�85�n]�2ė��?td�Z^dl�jD���Cf�}!P�nZ�Zsٕ׌����M�M�^2�%^Ee}_�ۏ��	aJ6��)Gj�u6��	�y���t�~�$�L�F��A �*���Iq���Y�ӕ�d�A) ��ZU�I����мO������[�u��
�]�ґJ,���#���R���]_܁������s%z�� ��X�4PDu�k���q�h!z�Nʜy�~���ў�-��X�H2�3ܽ8Q�y@�eY(�p����*����!����ū�)f�Mj���/�a0Do�םl+�>��>��Ĥ�k�)zz'�
|��5נ`�Hn;�;�mPBBv��t;O�K;0D��]�&'>��pGZo�-�T�G���x��s��<��%� �ɾ�]�)z��L�ը-��׶'gU�L$��fǹ���"b�vT^�����^5h5���!��*a �<�3x�W{|�~
�E����:E�^E��u��I�L��6����TP��b��O��a�4��G)m��pgU[��Y�2�)BW�������%t�
���-"�,,dԕ�sNi��()��$�
y�1�|�3�Wě$$���z����1��
j=A؂�Vݶ��:��f���AL��T	�<X�Z��pd
��u_��S�JjݪCe	��n�~B�U�_sc�
�ҟLج��%]�cS�f�鶠B��bv�4|�0��~y]�c���GhA����n(�:&�p��3��(���<lܨ��ȾK��Q�(�V�E|Y0��P�*���#D��E��'�BH�1�uڲ
�|n���ذP�CN��r#h�[oc�,��Gq�	[��A���Nb?B��`�ʔ���1.���3&�C~x�'�(I��i�iV{�Du���.���Lo��ɨ�xg�O>�-��,d
Ш�Ck9������&p�-DߌmG"ACv�U��r�O�Q���!���q�c�y]���U;�Q��isOA���`�1_�~�G�&��m>���<�מ��\"�0+�I���|�o��_{_���t��f�����cҎ��[�BB�lJ�ȉv��z�M���?��g�q����&�l�G��*y����/�g����� �����rc�u�f̳���<�^I�TMy��M�'��ܜw�奛X���]�f�="1���)��e/E������A/`��%���@���35�8�M�(v��u�����g����M����D���1��k��LKm0>����?�S�[��|1��L˳���O� L�Y=.T�L��m��p�lm��j��=��!�w0LL7 �Ur�1�<��J�X�|5%���HhYğ�������H&IեG{êx�߲A)(�-nqt2�3��Y�-ka���쏲�(zt�����7$��W���q�j*�&=��}y��x��VC��7��pF�Y8��J��i�.�����z/�v�g�
��V�����/�����a�e_z�F� �L�
;�n-
 ^X��WҾ�S��z���/^np�JEo��� L�]+ :8�{�4��Ƚ��6���İx&`uc
+CK����λ���O�GV�g<�a>=y�x��^N��_���BA�j��[�E��u�j�`��X��� �nV����������SRi���,��{5�_������/�D!i�q�56�S��������b�
e�/��`�����9X?�>7���(	����\��p�dy_	��ӭ�н^w�?Æa�O|�����}'��UC%X��:1%�셭樁�D�в������;��QyX_�7R+�& �����W��.��dN���l�E�V��K��@P����v���+W�4�nDv+�B�P�nd���;�~�b��a���:}�
G��Y ?�S<�Ɯ؛�\��EK�Ih���a��yt�],����%�Kd�Rs7������M5^Ŵ�f�����ﴩN_���(��^�<�W[�2�@���������-�{.�d'T͡_������Ks����}���3�#��Z��6N��_LC��byz�W������`ຎU<
���x6N�ϋ��Ȇ�9Ab=جE#�y�Zw��+��r!f�'��N˼���#�a�l�뻕��x��/� ��'�{R�HνAro����n�-��Zu�i�M���ҏ�/ �����+�7P=>)\�}��o��6C�[�g�a�l����,�,�i��9�q�C>[5��W)Xr����ٚ��?ָ�e[���,]~D`�e?'���+�^횘�*��h��Hf�T�q",�3�b�^��n)�A�rO,�����=�3���D~�D�J�Ͱ�3�
�S�F �AmWa���C���zX���3IHw�g���g����03oO�ڲ$\�Rhr���ۘ�(`�=v�E� �k��fX�{V�T�*�KwmK����H�G�B�~[����� �Ʈ�Cvn�	8B8���zo�1�Z��}4:�>b#H���8�͜e[���9P����;/�J�x���ӷn���Bv >�b�g������ܵ7��U�۝�� u�s��Q�lC	��� � QW��kJ�[�<fװ��U���h�@B��w7�&�-���S�9���/����+�=�,���;/�����LW@����/�r�Z�ah��uZic��BN�����4K[81'麅�Ya�_�+��kq ?1T�S�Δߗ�̾=N;��[���Yb��]�	7K-Vip$6�C��.�삭�w4Ѝp4�4�������E�������+L�1�ĉ�=���x1��H��� y� �p����u���Iم��$
�0�΍�X�4���h\�?�J٨�_�b���*{�P�*�m�`�d�N���/ ��h���_ױud7'�T��-J�Y�{w�+}ʈ����� (���*9Ι�GS;���sc.��>�/�mTB=� ���5E:{�
J�\�C�ް.m�'��K% �l���U�Z�5�r���ت5��-e�
T̨;�_I�7o�AM��S��xЪ<]�*ޫ�~��4����D7mv�1����KOA�y����YU��\�%h6q�\���j�`����zn3�mv�� @��V묪v�`q�F%�c��
f�Z�G5Z�,��5N���v"4�?^��� �~$�9��{D��3�䒆Ԗ�)�1��p���/_�V�踻�h������T���4*61�/\���^��$"�y���fG�ߔ���ɕ䪬hG�e��4�2�1:�j���zаN"��� �Ɠ4��#�%:o����)Nsc"��Y��E��_h�s�v��Y0�H�a=S�����	z���Uz����E���pb}��ѰO��l���l./'
K������w����W�w��J4Tt2pi �2��f\�0��߼*���KY*fw(�g�K���\����I�_NO����M�`Й�W�F���&f�	k7���3ӂb@�b��1�)����0��6S�S��G��Gv����#���x ����E�A�j�:����R䓟�d���m|�\�_���A�9�>�^/}%��Z  w�ƞ�"�����R�3��\.��A@1�g�J/��{���uXX�o'g�^T�Ղ�Q'�a^*�*T$�X"{�|xl^��a\Ň����u�e�J!�#Y���(8�&mܴ�4ڼ3�J����=���h�����I�-���m���f��[�Ɛ�)*� ��9�����K�C����������s�+���'�3#g��]3O��"�&=�o��w_j]QYW]����:0� 3Ü�i6���H�l��q�d�#%{��>��a��)N��s/��?r����bXB�R��8R���76��[�ɺǟĨB��DQ����RM�ѵ:����C�� 5W���K�dF y.9�X�B֕6+���;3�c��  �J2V�tj�WM�;F����g�G��A(�~��P�ųM2�`^2�ϸ�L`�8	�gng�D_�^v�j��|�2Z�  v o���V�9#^��T�3u1��V�at�0�v`6}���N:�Z1z�5w�t�J뿈�qJ܌&�b����<r?�8�ְM�f9&���P���?���Ӗn��c�_s}$l�[Yi���z�Vg�m�y�+�p����5�|9�٣��W�n��T�!�Iy[�]��Sl��Van�L�`_�^E^�]3���-�Ŕ��b��F)� pM�$�#��V��7�d�Z���%��V��6$ ��Fn��연rn��.�m��]_�e2��(��"�^�4.���0� �AɲF܈��\�\\r�M�q�ߩ���h�J���]�x&��AC�0��MQ.���i�6,�hSޘV'aWL_xW���6�2��$�����`rY6�$���&�3���V����,rX �����sV
������KݿmZ��l[��\�leHN�]�XA���/��Wwr;�#�� ���J6sG+]G>.�z�������4(1�x��(���y�x�T��K�M`=vm9�G/g
d�~��[�5r�E/[��W���ĝ��Ҷk.�����t�ߧ��A-��@�(RM�[��q���&� AZ�*�$0�[��ˋ\��	��~��ò8݇��G�2��*�)���C�)�����7��-�Ҋ��P�����*����-2p��!��ץo_㈢W.��(|wIҨyٳb`����� �cl�R(e�����Ru�/(^ϱ��F�i�#k�4$��B1��(�L��+��{%3�_!���!��sU�x/���j�N��֮ZV(�m�p��"�� ����������ؒ�� �J;`:W|75�@���c�C	1G6����F�mN��&� �5U�����l�!(t�"J��t����~bز�^fK�bgc��ҁ�F;��>�=Ry��BBЩ:	���amzY�\^�XD��<6�F����/E3`}�ٞq+v/���=�fD�s������V��7��Z{j9��%�����e��I%X��[� ���t��=3�8a{�.x�R����K�j��H�m���}ʫ`"�ڷ�ђ�N��RV�e�A���z|(�䴫����,�9)Amba\i�$b��|kJky�6��VK������	/<R@;sV������6�[8�!�H"���%�)UőJב�^�4�oJV�hǞrO�ȟ���p�D�+�b6u��e�x���r!Le��w-�1�����'����`���SLS�
Ex��R{ �('j�}G��hn���
2�BU��"9E�M���3�z�^ʵ��? ;0�	7R��H�X��H�h���C�`/ӂӲ2;���p]��pӰ3�Qt�CP��9����^��L�b�!�ŋ* nb�A�����&��ɼ^�4}=�Ķ��%�0T�y"�c� .�d����b����-���Z���Ji	�ưE��-��K�弌95\�NXWFG�Q���b]��}��c�"~A��/Lʒi( �<r0*�ǀ�W����x��v\F���`|"�,�O�1\A�V?�{	]�+X��"���[���=�p��	;*(g�%.̹�]?@�C�ǳ����N��	gHB�<���O�Ll�b>1���Z]� �!1l��DlP�n��
��1wNŘ�SZ9�Ccl�+�l~�ˤa~e�%�H��OЕ����fe�Ϫ��	z��1��K�����[���2�*�{�G���ɭQ^�|�b�A�L,�]d/4�P��� �q��p��s��B=�2���h]HM�j "x��S�I�c�!|��7mu�<�K���GzC�l��3�V>�`�\	�p����v������V�n���1��<�e��Meg�m'�m<�__���Kqˢ
KM��
_��ru�˃�:5���Q@Ѱ{�D+�yC��!GEB���{��|%���եK.�%��:���M�i��	�Ymp��u���M�Y������v;-��[~x	�����9��q�N�7�l^B�Y{H��}~/^�F��Q�x��|���65�XW����T8��6�Oz��E�⠍��xˁ���e������1N�/t�Eh< k?64�������\N<5�D�����@,6��)�`U�SSY:�`��E�	"���Ty~e�q%�^(m���i�3,���e��0g��G�h���Nު�$����p����
?@a�٧F�?��~��8|(hQ�����������nxUm	�Őf�v�f7
�x�X
 ��Ū�%�A{Aұ��n��L3���0
�m�Dc�E��L���Q�k<A�L��<�oV��F8U�p�	�C��*�Ք[p
�^��d�E�K�?�����v�b⑇��Q�W���2����eʣ���խ~!y�Um�>z�b9jۤ�����O[d�;����X*�|�A-�z�$�05��7�ԓ�J�6�����ϚŰ���A_j_t2�3�h�Cx�}1�y�q��a��~�4�=e��ݢ�6ܐ����J!t-��b�DC!�T+���o�F�ʶ���v�_�5�w�����l��o��� ̾|��sB�t��]�f�)�^8�.��C�)��~8H?�C��/��7���`;��GT��O�h?�O�(lcʕ.v��TB	�Y� �i�"����2��+w=��?������>���Z	���K��TM���ջ�kV��@��(3y�0\������`��jg�f��.X&�q?�!�u�8��׋$&7�"��;~�� *qh�Ǥym(��3q�%����6��;22�tޒ�a��������POk�NLધt�}�A�v��q�"=(:�)Vun?7�P�q
<�jY�O��2���p�N*ON��!�]�3��&��������胒�q�⯖�2+�pH�DiW2�����ю���Zw+~�Q6�t䥴�@���X�l�֣�4�{�w�S��A^�ů�f)2iI��R� �d�+L��K�8��N3c"�z�R�+޸4+%ۈv�nlR��G@/�@J��G!�4���>V�si�ȩ�T�҉l[׼�:�2��4i���c�XV�B��'�m��3
�oO��b!���ݕ�5�Р��O���5|u���p�3"��Rz�(D�@yŐ��R�]��b��y6$�%�Y0�\;�
��{(=M���fh'g']]Qc�>S�u�{���������|5*𥔛j��/�����,zҹ��vC�qn�+������R��w꺱�Xs�n>���rO�m6�ު)v�56ะ����������Q�I�G�����+��-|����@�b��N,��G.�ŧE���
j"��.�x��v%�nX���x�2QB���$�@4�F�H�D^ف.ׯ�v�h`�������51}�H��ۘ(m'�����:��j��R��-}��8�����>��[����Oz�$�V�/;)���n29�V-��"B�|�I�Ӧe�zy��XC��iy�*��Z�"i8�=���c�nŞ�	�AI쮇�������Q>o�E�j(;@9�++Gl��^�};唿��$<u%���>Is��"��ųY��k�ax,��f/s;_RK�S�6������_���������0}�:X���u/�\�`f���6�'\	�`�m��9s�Tx����Rw^d���O��S�������5�^+��SV�=`_>��S�a�6%J���X�G�Qc-s��~���铍�:T�f��Z�2:����l�9�k/N�LZ������p�d�욾�bX,T�Y�>[�y�jE�!e{���ܰ���a���ģ��)�\��s]w?�p�!Y�E1$<�㾇�"�F����<��׻Ȣ#��N 4~�{Ã_��Ȗ�����Ɛ��t�+�@jjG�= 8��~"��^Ho��s�?i��S�}B%���8�9��}�6R�ē��}3���n�!Q|z{����b�0����X���~�2�'����{O�cr� u��AM;��!R�D��`dԔy�t���p�:�~�����O���JQ����B�u�^sx��FQՊG��P�� [{���R+��O%��*|@q�$?��o�>��Fb[�H��T�Ź��]V�Q���^̔���:��Y�"�2�--��ӊ3y���K�}�m�B���� &@q�#"�TK���>��1����yks�:i��Ls4�Z�jɭ՞��c�a�֤�n�x߷:3v�bЀl�<�1;�A�Koi#��B����6�N-㫞���k,j>s~��L��h6���V�����; J�=A�bl.���s�wE:�q8���M���������S��}֋[02ϐ�XY���0Q2���((�r��W�C� 3���`�i�  DK�3N�����m#s�����H5�;A-��SS!�io^<r�y�5�>F�xz���)܆�'���n:N��j���X��zĎT�?g�C-උ]��3+����3�ھ��>%���)���1�9z]�(�ۢz6��b���Y��*�:���ح@HI�qv��%{��������y-�fEج�|B� �P�@��w��q��	�2c#wxk+5j�N�{��t�ݒ�EEu�j�B�s�s7�'����fpv�������.�|��f��
+4��K{��'Tɨ��q��\���0�>�L��e�p�C��5\P�A�)@P`��Zk�*��gFD���\7�mb��/�UV�:�|�^Ǒ�D�\�e�7�H�}y^Ty�E3�����k��ǯ��y���x���<���ɠ�1�)�SC�م��/2��f�'n�������d�F�+=��$���S�eT/���rA3$��I��=g�vV��̝�A��`���M�<�����_����bu%[�����lp��Zˍ��qh|;[<_X�8;סB��Mk(6�C�4V������ڔXiR��d��~��p�S]v�n��؁���͔���mR�X����c�ZC��m� �4��ˡmI]hL�a�,M6@GS���Tu@�k���(k�Cq~�H�M�{�"��ko0���1�|RLzWH.�82X��w�n�w�i��CZ73���\Y���jC�;���=T} ��r��6��"���r+�W@el��-�37�9�I�@U�Иm��ƨ+4�{���spL���?|w��Hok���H�rA@^�Y��z�W���8��=�Zd:|��M&P����j�C�t��8��%&_�'�,�p�क���š���4�6�s���yA���n��v�A)���]����QG9x�E����_ر�]&�"4�RVkUav23ܘ�X��c���3X��q g�}�;�ن{22L�P��FGo�ˑ^U�/i6�N�i){Pqk�N>q+0��,���G� ��gm�R TV�X��ղ9��k����zf7�e�HAIG���*��fN�z������N�N��|��J�ϲ�?q{��y}�eK@z	�	�p�6�A\̴w�wL���n�1c�'��>G��2(okN�l,7䧿��r���q����w���T��r���[`D�mwj.��5}ݗ���9zi�ly�M!�������;�W\��K�B���s��v�1j�M�CE��q�x����<���CSJ��\S��	�i�WOXgu|�`s� ��:ųX��uXF"�J������h7����0Q���>��^�w���q=���ec˟��h���BFcO���ۼ���r�����]9�_�:�gb`�kփ�"��7zGn_�ۋ��hQ�k�l C��o�q;T:@��/{ɝ��� 6=B^���r��{�x ���mA��?b�I]�G�[��!V\\K}�~�8� 1;�O!��p���Uȧ}��� �&px>�o*�t��G��߲���mB�������!����
�sֽ�`:VM�*4x�6�o���.���X�VN���:�����LxGC7�G�7sF:4]el(�U]K# _=��z[�2}�O�zU{+��b\_�Hi'
kL6��:�C?X Gj��Q�t�L��#q��"%�b�Gf�"1{O)��ni.���_ѭLu�5��j�U`tkL���`��R���$��W��sk�:{�����c��v�㗷#s�Gx_�)�W^=%8+c3�K��w�H��oa�p�X��55�U9<�Y���	�_Y��!���m��o�UDO363�F���p�f`��B�i�]6�_0��J~
�Q����=*���9J�gf�yz"�1�3�o���t���9�W8e���(5P�3�}vἓ��lE�U�C�����9���n�u��G�L5�CO�գ�Ԧg�e���3��
g4|v�M�?�a鱔h'�����g��y*�ʬ?�5\MԽ���ĭ�����Dт��+V�$5���-@/ͶD�܌m���"��wg@��F�G#Ǩ����?}1;�	�����%Ӑ�~��+u9��<
T	i>'���d�xq�)݁kz���<��|�[��?/k���cFay�R�����bX=��&85m���x�MЎ�Nm��2��*���}%�L�թ>xfyNx_-?��\A��Y*�fJ|h�spP@�& d�k>.�����t܋�uT��M�mt�I�1����	�8��N恆hA��y>�Tr�Pz�7���2\�_ǃHrZ�s�>�T���
�
v�D��!5r��)m����TI{Jߘϊ���H�ؽЃ�yn�2�6?��4;D����L��8�дV�W ���'�� ���\`�����4����l��d[�DIN����jC���c��Z��Dx���]X*�G�W<��D�IsR"b\҇�����`�N��H�������=𭤎
xz�%PD<?X��]tqM��u�ٔ��.��"���P��-�(�ZF+���g#�\�3��yb� IS{��;����J�M���9�d��>E��|�h+�f�(M����u�td/!�a �� 7Rr}sCh�xݺ�,͞�=%q68��Y��/m��/�pa�*_w��ʧ��7���heᮉЏ%f�>��Sy��B����5O���BH�8{��J
 ���4I�v|��j]�{�cGV��n�KW�*ǂ����! ��@��V�;����3M�g��e��Si󅖏�͍R���4oM��7@j /��S[Q'�?2 ���qr��\�;��^��^_g8K�A#��U�_���([=�ߪL���g﷼>q&à/�I������j�n�ƿpN�ɘ��b#c�6!x;9YNl��jӼ��T��;�����9(a�)TV�i���1仟��� U��K5I.P'/+�H#���S~����PՈ6�Y��Z�
��G�t7�T:�^�R����,�sAu��Ќt3|t1� z�i_H�鐶�
D�}̈_Ae�u�t/κ��L;��w��r�<�P�{�>��eB���ŋ�q���+�y���u(���P�e�Ƞk&a�o��?�ag���ba	q^�g���ժ�R�^��Ԭa#ﮄ����p�\�AM��g��F/r��~��)ak�4�q#Z�?9b��\�_!�@�[�=?ܶ\�e���+���������Z��l�>�5Դ�#�T��u��@�z�'n)Ȉ�t![ t��NQ�O~Pt���g�Z֑ו|`9J`��in��K�(d�P=�$�	0�"D�z�a �� >^xW|�k�Z�Ȧ���141*4Y�r�����8��?�pR�����R�T1�t�O4-�>�};[Ր��idm
>Af}X���,�1�-9.�[���(���tK'kU�W*�U��I��>���1K9��N��*:���F�����_'(|�Mvz[c��[�Ao�{�"G�W�����>���[�0��Ԫͷ�,3�a�.0={��{�k� 	\���V�`���l�̲%�H%̆-��2$�����lW���#�`����I��d��C��VmѐF>����QG�:�tшq|���>PH��J>��	� ���F�*��[Tӟ��,��Zf�1�tJOE?k�Ћ<WI�5�����n)K���S�+ܩ��p��[���pD G= ���ҳ(櫼���[qy� � ���H.&I�k�h#q�=��Ǳ��?�N�![��"�B���j��8n�Ȳ *�kRd��n�%Az�Lb(t�]J�3��@�����!IA�|�S&�B��/P����${g�'�Z�Ds��NB���\i��߹�Ī��-���/�;�nAZͬ��b��]>���3HXa���Op�!���g�a`<R���P�=���EL����
sO)�vO���}CVC�GE�au~Js��!Z�|�r=�+'��o)��s[*LL���>Hf�ZwSH�Knܠ�.N��𐱋��OY8��gQE't6��V+0��vc[���D�����<�'l� _7��g�p�N��Q#�4H���U��v0��j[�����¾m��tM��.U�Byu7�2@���f�me0���,6I(�q�z����۪��5�T:EvZ0]vA�/!�S�]aC~����9��)��5=�(�� �	���.�Hlh�,[�V~�j6'y�������F}�	��ԏw����a�8)u&u_��$آ�>�s���vD����9?�l��I��m/��\��;1/�w�BZ(-��\��+u���	��N�I����p��ܮ���^r\'@B�I<-a.����As�F��(WG4��I����d�<�T�@�����o�z<�m���c�G_/������;��r��y&K���=I����1kF-���v�^i��J&�-lD���s�����DM�@rd�>�Uz�5���7l�6�7����jD���6|^d:d��M��!Y5���:��q�R�˕s��c�-<���n!d�����\�4��;��P��sCPc��Z.�(ɒV����3f�"Nmƌ�iPiT{�Ge����$���[�N�zQ�\sY=���c�����=}:Q��ܢ���)d�M��F��wrEE���d;�z�;�����_4�w�Y��!؇tv�Xm�y�y�|���G<���oP3�n��վ��yC���W���_�L�W�����N�ef�4��A��y�� �җ>�oV��3+�È$ˈ�H%I��J��9nN\b���(9qYR�-v:�^��R�#(7S�Sx������M��b\n�!|6���=G��54�Q����ט���v��Bv't�f�NR۸7�Od$��q�1Kb���h���G��:�t�ʮ2� �ۘ�&�'+��V��'��K���B��~�&�C��r j������ˑl_��_�aQ5O��&ZÌ Ļ�R�6�V˵�h)W�c�A�O�	�$4j��dGY�2�X�?��u�D���V��S6��z�U<
Ay,�t�*�MiQ&��e{ @���D��:�w|���x�c�(s�_���$%��<$P[M�����˛Hڞ
�Y+�_��Q���c��Z�����s���?�5��S�VT	�4Pz�� P���z:���OF*�a�W����dCv��f�{���G�9�Wm�&�Y��ς�}���_��J���6&x�g|������14��,}�?�@6&[�|��O��ҏ��~�2CGtᴏS~P;�$�^��m�Tuu�*L�X��J�NHvJ,��n�Pl3 ��ɻ���&��6m�F��� n\6�8�����l����Y�؆I�ߡ��nQ�$gwrْ>�vG
1�}e&)ת]�*Q7��,9q1Q�'˜�B\J�jI� �R`�a\ܥ��mP��׊%b�ϟ��/��6�^�!�࿢�Om�Z�g�D��ߟ�^sďW&%��ŉ+|	����".�L�D�W�p�L�B_���9��{�H��X����Sf09(L8�q4�%���p�d�΃�LDrA��������y`�:�^'�&�1���k.����ϟkJ����ee��?�%�'��0�D�k<���B󼝈Z�zW�ˠC�!�;�-��d8�<(���b��v,���׳+!\��rƫ����S��
�������5b+����꟣?u'`�^�3�h�5C�J�Ua�-�uq�as�}ITI")Co��VH��j+o��>.�{Jt��v,rh'��NGN�v7vx���8B9u�Cȕ#�u���������-eSk=tF�~�6�'�Z��`}���=~�+�7Q�N2J�w�}hĦ�,H�8�M�]�!̶�ѤF�*�qO$k�o�3#z��1I��5<J�Q�Jl�f�aH����pq$�Ð{<z�9�/���C����ҝ�C�iN_���3��u��a?��ꅸ���'?iw�^6��l�uX���_���(ڈ�*ڛ�O[�����a�c���9ӅO���Cg��%stsk�5�xc
o�5�]�D+;k9���$�+�9S�R.��R�ր}��X?E?!�{S��.B)�3f`_��|xO-�nd�����X9�ٿ@��쀫�WX����%:)���r*���)���oV�����~2�|~��f2_mV��v�� )F�!���V���sa����,Co��c�7�_��N:x��/l������0�#�2�
��D6��>�f%���b��i��Y=-�W�oi2�v?��Z��1*^�y1�]ŗ�^�>7x�BL�/U-ǽ
�����cF����� ����zY�v��2M��Z�i�tMr��ϻ(T:��Ę˓�8!���ٚw(=/ϹN����Ī����v�'�lB	&����(<Pn��T+���/> �� ;��ڭ��Va@�E�������3��vhSx8�w��o����!�b�4�uY������`����zx�fr�u����h�P��y�~H�a(3�^��G�?r�\�Lc�gK���L�2�q����֐9`�傝���*	ؤ�|�+�h����M���*W��o#XA�3��
bc=q-k�wJ�׈]DIC�,����%2u��#oNxQ>s�}���~�����t/S�x��aJ�l���
�7t�z;�a�9�j�4]༢di��[�T|//lƦ�5~i�����_i�Z�47Hx��0;����#&����,tK����������®d��i���8�72�/L�1�L��o��C1A�v��׸g��B�q�b!��� ���SW���{�T�����N�.[�3C��[Q�B�.n����Y���
�
�����=z���H��^�0A����ҵ��"m��(a�
�uڛ����� Nʾ/T�D�Cg�I9V�`�{�dg��m�Cۃ� �}n5������3}~+1=�$R,pcl$�H<��_	�*�vN�)?��	S�ـ�$�V�\�G�0�gOJ��z%A��q���;���.}x�J�5�z��.�A���[��V���7=A��O�
%J��ͨo�xͮ������=�Q�ku}����fZܝ����G�V�&����=\�A�� Be�tR�q.l�^+a@]\�3M;���ڤ��|=ƌ�<F�ePҮ_�IU�C��/��}o5f�CNl!�`���MuWҮ�dsy�J�X½�&�Y9�:�1 m�k�s�) ��UH��N)&���,���A��`�G�&�=��q�K�dPQHMf�7�)G�*#��꽍7:l$jbL�i�㦊���	 P���6A��`���}���zg�4"�&k9���-���3e�iO<TI7�3����Y�����g<�qOS���Ne���0s?C�-�SD�����\.`)�������:��ֆ�.CɈ�לԎ�a? }EX~��I�i�w��ӿ�G3-�s�黊+a\rj5�.���nO<�+�OT���]��teӱR�Z�gF�ٺrL�xH��~J)�%�rg�3���?��7���;�@�(]p��BJ���X�_�/�O�Z>�#I�;��=�iUs�q-�r3�\W����-^�Z�UdY���ʦ9Ϣ���v��y�3X���/>�:�8V��x2����x���I�;_�^�E�G\}����aq�����\t���^7��������A���A�_e�7�C
�W��XΝ�yR� a}J�jFS�����61?�N�8b�H�+rD�?�!�E�5��<v��u�r�yZ!��	M��T�)0��u�#�a{�\T�%Lz��FE��=�o����Z��co=��.�<��/H�a}���K����I�б��&�\!��ɝRe��ש�&d4�)s�-�w���|�v�� �:$����u��yc��$;▛K$K��KU�$pԽ�mG��kc&��!���X�2�}���Q���ᖶ�����@��C=�ŗG��)fب1	ѣ��%cdo!�����bP1�RS�AU�1-���Ӝ�@�%5Z�E�����Щ���0��xT����\\�����>?�qǿ~R7� cV��^�HϾ�����z�
��ʍQ�K�	�$o"2� HOM�Y(*${�]�}qL���(�(�]n�����W���~�Hz�����I��f��yZ���������ICY�i]+�eh'N�..m'|S��B��#%��g!J��O�˫�f�O�`�����;K��%T�]8Yw^��]z�Ĭ�wrBI����tmd�q���jb�{,��v��t�2�8>��eE>�ZJH�`c0����.��ܧǵ���%��G-��*���w�ʟ���[�e��3�>zhV7����� �衻m�m�hQ�xm���dݭ�r�7k*��'�N�7�-y����a�-���"��<�e��fҭ�3�v���	1�(�殦hϯI3;oD�(z��pf��m�����ݤ���nj:,L�!���T1kYT�123��ێ���T6Dc��#
���9B�t�	�C��/z��ك�G���핊`���ia�l䫎UMs�*�tD=!#7�&���������D-�rt�&=3��[˩�m�h�;S,^2�[#L�P< ��FZ�"tm�j���W"�'rBz�-�N�:I�r8�\�P���BXr�U(1�q����s]�׻�	Q�VL�ܠ�5�U <�����a�x��W��DY�
�Y��ը�����΄�L�p�ޛ㗵���(�D��������[V΢;��`�O�1�v��l��Z%b�v�ݾ���:���f���-�'�����]���)<P��&����,mJ�@�h�Y>��ˁf��������	#�a�RՎ�+�������|������*�p�<:c$k��O$<�=�T�ޗ��23��͗JI��/�P��H����RR�~ë��M|�͇�$Uf^�Ϫ�E:�/G4>��Qf�Da៣7.�HR�z�RΟ�}�~���x)���i	
(B�Ol���Y�X���$�R��Z��eΥ�]Оu:8z�Ӿ~9#�������!{`�AƸI�_�n�ڷ p��f�v�鲬\	~'��
�t3�S"FDe'0 Qs	�FU%�7�v1ٓ�@�-�s�a��sE-"�v��Wpdp��C��,@O�n�*v���I��0&MM˛%h5�I�r{4��9�k-����K���xiB*5��l�)K��	��m&�ZV�x�剩{q����v��a�怍�x�8/�Ybہ,���>�_>�a����M/�fJx!� �U�,�!\���3u��6�T�~$��F��[:�F(���e��Jm.���7��F3�!$���<ȿ*�QI��Z|0+�����D�Ò8^��K VS:�����J���~y@QPP�Q�|�~�V��/'���Ƹ��w��j��y_&}�k���I��iA�#�A�C�ot��%���;M(�v>.��Yn����Y�31�������������O���Y:�A�(���6[FB�b.�v�m����iE����G��	l�ag�^�h�yu��l*vx�ߤ&�Gm�S׹�WAݟ���u�z�k;���g�
����-)�Xe����e��	�XdW��h�%w���%�%��vC�A\k�� ��f�����7����9�Vtؒ'�5ŨN��%��iAO����=,�6f"�S�����Mد�n�)Z��P�ӊ�����
f��B�di��=���F%��}|m�}n|q��]��ʨ�����ԅU��f�ߡM���leT�����v(�7-���d����y߅?Q��,��wI�e�	ӱ8"#ݯ���{VJ�}Z�h3"�^&?�F�;؈��:&��එ	b��j��ٷJ��ܬ���Jde�����:]�(}s���!�wi|9��Z#���Dca�q�Թ��J_��b	U�,�a�����^�1"��}��l��|��m�l���j��$ך�������L�Vݧ��no	��.�}
�f4���%Z᱓�⮚ɴה�o�K��w�oYE8#V`�}�u�����'J�oP��z�݌v��OC*'NBS!y𕫏	*9��ґL��M7����_�^�&Y���n:���IbM6n�F[[����pn�^�t-O/$3��.*uD��Յ��mJ1��I�0�����	:�]�Z�0����e��FiuN(⪭��77Y��ӤJ�h�Y�/M�#�[�k ���k��&����q��Χ��ξIX77�R�{�Bp���v`��n���h0ܕ��.��P��BCֳ�㧤є0�3�%�T]�4�����nY����9T��n3���82Ǯ���t��X
G���Q��V�{N벡�mn��\g�j�-�`�m�I#��~"�}iv���&L�G0�'�(ة��S ̖Ϋ�T���Ӱ����&���t���gc� �\P/�{����m����aτ����3V��8��`�����M��u|�sZ�k���F��DXI��{KG�3�ͱ�䑔���������x���E0�{#a9G(�Uy��Xg���S��2�+h��
݈���J
�@Z��
=mټ-'��u�4�Q�źt�lS���אѳ��vZ���s��f�zP} �1�1�)\?������6�c�/�۟W9�@�����m
٦(�ʶ'��>�A��R,\���^�C=�6k��tz�9��;�@e��t�Տ�ȹ�܁'���t �w��Yt��s��=�g�~Ӵ��������� v��lz�~'��;�������MFE��_��Y������V�+�|�b�ը��BZ��������'`;P���<��5��#�1�p�>�Yhyo��(���ی�UppM�䪨z��-x��w�3x��OŬea�+vgj�'*>"8m�1֗/��M���Ϳ�$�ǹ�A��rd�����)Ѣ��	����c�������˚�.XB������޳�*m	2�{YEέ���Wf�̳�Y�GI0��	�}xS�VO'y�����'2��W��``�@Q���%[Ve5�J���mzg�vM�FΏ�H(H*asW9��Z�h�@����Zn�R��3�(I����_`��PD햜�Ґ�U�{���W�#��VH�����;JSn����=��{� W��~������)��)*.4�D�)J��]Ja&��|N�@0�L7�PH��	�oRn��'������w����<OS�Yk��s)�+�$%�Kv)dE�@ �H����wQkPz2p�R��Ư���
���V��mHچH���+��y�Xy�V-W܇E�pՋ��i��xX�w�(���qa�g���c+�i]��O����tؕ��=��/c�^�´���X"6K ��&pA�����Zٺ�z8�*�B����s����s� ��'�`�
��R�g-`�X�=�:�=�>�aP��I����E�f��J��̣�RLkz]�&#k�+���i��φ���;�z>�Ԣ��7Tz0c�}��y��gPV�����:���@x`Ns��O&|@%6�� �S��g�o~�M"��Ϸ�%����Kcc�@?�2Y�#XZ���xF�S�����O�7w�o����T먀e��D���L1yV��(�G��&J5��X?�1��p�H��q	�'T?�Ėi����2r���U@���#8R�m�[q)횕��Id����}B6_A�0��^�=��ep�����*1u�;[���(8��#(IL�i�y(�������"v��M�ꘜ���0���w+�R���2����_NQ�H�+E�u ���yW���X�>
����=���e6�U�ooK�-�W��ղ��&�p��b��;�@����������6}��Jyt�t�pOa?�I�K��#P�n�:�FV����L�1�f7�[	o�B��`�4��/�q�EK5��}�T4�
e�͉�����'��d%,����ے��'6r"8��xD z�jߎ����H�����|�X�OEYð�Y�k-[�d���-T�\��I�S46?is$�Ж1Ʒ^;��α�r��DbQ8	����"��׾GĀF����ݞ�!�Z�$(,۰�<��5�?��,�Ľ���� �t�)��Ӥ����4f�a������,sw��bu�B�c�!���W�^#���t��:$��^�]I*�}��\�M��S|���P�V���OZ��|MFu�.�P:GW��
䢣o8��`��Zf��"s#8˦�o�ȫ,�TYF��&��l�f�j_v�A��5\�
���U��l��e� ��3.�g
������nr
���T���0������tnܖ `O.Z3r|�L�s�d����1�w�9Ikt"��z����G��������^�����Ż��0��^�"N��6�~�)/[���H��Q�\���W&�ÜJ��>��l���CO&O)���A��A*EA�D�
,��Q�6̱|�,{U;V���z�	�V΄�/tn�b��+�X� k�h:/.�S��֜�nR�J_=�)	�8a9�å6I���ǆ�MK��A�����K%��0�*Aآp�63T���"�2��Y^�5���0,Tڀ�^���B����s|���wi���D��l@��CG+B�7)6LvXS�z�'�����i���;]���U5z+w��?�Z����iz�kb2
������fڀ�L�~&��c�a�%���8ޅA_A����mm6RX)�=4V�X��%p�ZCX�l����z��9���}[C��Y5L�T!�ӑ�va�V"�k!�rTҰs;LѦA�\[;�9����?T��t�b���n��9
;B����J����Ֆ���d^첾�Ŏ��������(���\2��C�	0�ynad&�n�b��m���L�i�K[ J9�[0��Q����?�"5�+C�w<���g'��faHX�E��U�M�٪���\�2� [yÙ��s�L̔QsB�eE$Ly���l�Ҭ0�2�[U�5����I�t���;R���.�;n3�A���� i` ~�O��ǌ�+�Z%k�
ٕ���
�8�hɿ��\ �#���I����(J)׭ͣ0�  ����[��a�V�E��}�B��f�X55�W�1u;��<M3��@���V������h@X4E�%�P�e�v?��khBDz�MJXUF��l�:rW�G �³���<���N�5tD�\g���u��yd�t��h��a��*�O�Y�IYS%�Ǉ҅w%��H\�����&ҭp�K�G� ��63
�}��}7v�|Սp�U���0g�0�2�uɻ����kw�^5�ꅴ8���RUμ\v�;��,Qv��X�F�V�d��.S�.oU��HG�S��������a{��%�ca�0��˱�R��f��,ͳ����Z�Ǻ�τ>iji?p�J/���f��@�wb��uZ�.�|!/�7_�B�ч��(��#� r{��U'�]��g=�2�� 2����+*��h���L~� �r_����;�?�&N�RDZ��A��m+��tkRx��^λ=��"���k9�'����UN�vFѯ^HrDu�!��R���隱�V���b��������&�a�q��i޸���hi*:pr���F��"��A�HؘBTׇ�ê���j�0�(��a���&��sգ��/鮓��ݠR[�~��]��I.���'~��D��ϳL}g��
Hv����]�'��������:i�v΄GE�ͨ.�bw�!�ue+@)]
�Z���M�2��2��<h�҈[K��Y�C)!�hR�	�Q_�T���=Yzw�S���yw��j���7���~����E6�ܣ��Iß�fw���A���Q2�;��[ �-��
{�s�}i[K8WI2;�1�C�����B�����v�+Qڎ�l���-&+
�a/�O�S�"�����#<{�zc��y	Q��x�;�&�ʉ*m��Mo��e7>����O۾Q���/���b_�9�ќr�E{����$ځ�5;В��F�SXŲ���r��s�[R��9U�Aë�Ara�h���Ĝ�����^�P�����,��<Ȧ�i��܀�R����:VSle 8����V-2���G(v�>/]��l��h�Y�fU��NDJ��?�V�����>�ޡ,�ϡ��C(�(�!7ͮ��+Og�!��GR\��q��bq��A����p�s@�qܻ���>9>j��CE3� )Kf��fo��<��>���i3���2�."����V�K������gG�kb ���1pz��j���~L#�8�dؑl�L�!�'F�1i���lokذ��GK~O��$���B�X���yy�bmɕ�b������[8Ts'7�����os�����l�M�x�iҶrL��O��3 5�@tc�Y�.h��\��:Yߙ[#���	T�:m8#�uĖm Y4�L?��H���V�	ؾ�Z2?�:r73�@���MÓñ"y�a�)��ρ8�M��.�Ym�I�ٹBP�p�u��f�;�|`G��l�������=��vK���iPs[Z�r&pq;XO�8�:�H�B�&Ph�j.;�A����g̪�`��~1y���/?��7_��e�b���?Piii�5�e?:�ù@/},�/���8��9��N�x�b5��u��v�5��[� U���U��,"X�I>�:W:�N}t�v�N�6H����y���R�W6�5K\3��m�#>�!�� Ė&f=�j: OA�$��;���B��*��#�#�E,�G�RV�o0���cs�U��Ć��^)��0�n�8���������jt ��}<Be��)�@�쀀�8X�΢������DX����D�O�^!R�PFd�.%"�H�if;�7H#X����m�n� CJ�ⱚ
� �Qc0�W���q������[ W������X'��oy��&mނ/�O�^�a��j$��H1m��H���)9+�I�.�D�p ���[Rt����|t�����T.���yJ�B�R��X0෱h ����r��s���ʾv�Dc>�8�?3�<�{����o���H�l�O΄��z�؆���K�\���`�78;�ݒ���?������1'�*�X�s��#��h����i@�{�%[���6��T ыRR?�����[�S�����f0N\
�#J���Q>c��)]��*k�u���蒍pA��r�+#?�O$�f�It*;�l^�ə�y�g��ݐ��V�`�<��<.>�f�*��8�	��)O<W2�p�榉w��
kW&��:ú8�?O7A�^7�����ǉ�̒�m���G9��sJ��/�>R��&&�N\M~�D�Wԩ�y<Z���:IĆTOv%(<�p�9k��A��2J�r�qL�y�l�< �鹢�{(f�ج���+M�����qC�ԽAs}Pbd������V^���[�-�7~�]��5T�!u�/�d�y��
	c��ꉼ������m�`�R�M_$��'E����,�\.�8 \eD0H�$o�;��pR	,���(P'YFy8�m)9u�'.� d�yIڊ�T��
�1���e-#��p�+�J.����L3� �?9ϒk:`j�{h
�C�WA���{�s�H.�,�R�=��uj셾]G���e��;i7�n���zV�J�H��w���sHw�3�䕸2e�'!e�<Ep�f�\)JR��n}r�����Ȭ_^Ӕ�ٱA3�q��^�$��@s�W]�Go�]Z�0�	��: ��z�t'���0qXZ/��5�;�I0�5>~��[M�\�e�2���xzt����eL��XFbS᫞��T�V*�@)�h�+��񆇁�5���WH�'{�?'%9A���FO�L��8bWP�"�	��ɂ��*TU��C˺	�)�˚P�C�V�#!Xe�����:�9U��*�z�#G���M�OÖ��Hb��a��.���#�)���SYAk��S���$�%6�ɍ�R;��#�񱪡�#�^:�]�7�ݱ�&S�8�_�=W��۵C��������Q��*xFo�Q�������S�*�k���~�F=v#9�S,�x��K�0RÞVxr�UC�m��Xq+���Q�u��K�А\���q�Ѿ�$+���j�6�'q?�,�a�{б�������{�1GV�a��?XB�V�6Q5J�B��mg�VHߪ0n���������f�Xc.Kĉ���\[1��.�v����P*����c����Q�,*������x��	p̂�҃g�Iy����#�?��F95"�$���W�墯j�iW�X@�^���F%�P�,�z�jq�'�P:һg�FB�B]���Z���l��]�����"��\ �<��f�j��q���������W� ��?�R���W�d�#?��"����U��}{Wݩ��~׮��P,����M�=��Imd0Z7��P�S�0Q��W�����~�~�e��R }�������"d6�*�Zww��W�o�p���f*j���r|����LҾf�|��C⥒��ITҴJ�"	���\����4�ӏ"��8�Bv������+��\�/h�܉e��L��B}�����jN���u�O\ Z��\�`
���N�`%���4��-b���Jf�n�J�f&������	��������R�U$A`Z�J�����g���Wc�%d?rΧu����u/���A���]s���`�\ƃO�R��"��N�-u<	S�J��������pL��q�� Wo�%
�h��F���'3�-Ǟ8h�o�_���I�˄�[Ѣ��D���\iT�Z����2�^�r`�㴨��&�b�{�
6X�h[�VR I	I���e�G $��
��.uhEk*�Wv,�J��1N^Ä�ׂ�y͙�UM-h�=Bm-!��sb`��h|�7x��ʥ�MR�o4���^���6VH���'����7J-�C[�R�}c��S�e
�p�i#~��E3/Z?M��X��9p�O�(՗�'���w�v{�Li��?�5��à���22��U0���(j߃�Mo������˪��4�N�Z�+���Q|�y�ˉ�^��!&��� ���'Y���RYɲ�Y�v��c����;;�6��_�D8� ��Z۝�L:��/{8J.v(O-�R�$���N`k��g=d����+.x[����_D�.1�9�;�m.ZҼ�θ��(���{oYCY�"F�:CO�N'��慌�F�,���atMJ�ģѵ [~!Zo����6*�v�Qb�p��5*�O��xN�����G�} �;� ��fU�や�Z��X�&ɟcW���ڵ[|���an{嗟l/�6��.��z-�����e�)✌��;l��[��]Z3T-tmE`[q� D�^6�и�K�CQ:�!t;(�����8٭�@����-�4I1@�UX��n�����j�@E��d�s�7w�P�R��A�5�Cl��x�5i�G�9���<�a&7H���O��o��h�-�Va*�A�R��i����eT+�!'#����Y �C��.:M���1��W�F�����Sb�nnc�`������d3s �I�:�!q��m�A�[�h�!uDwWB�V,���T�XCeU��(/u��-84)I8�z�M�h-���2ʾQ�0� l]q��(w���J(���M��\*y+P�9,�N6b���(g�sam��n.����ls���q�����Y$!�{�'a*_��mDĕ&�Y�
���	�����, ��XIe�r��E��v"ν�v��ǵ�&&*U,|�z��ת��Lm+J��6ϴ��Y�����A�֥�&PFΰ��N�|��r>(�� }`|c���<6�/_����B�vTo)����^/��s{�qJ�N;æ4[�e��$F�9ї�L$�M(ƌH�z@J� ���$��C��T�����B5����C�����׮�Ω�u�;��'�F�-�Gu\u�,8+%BP��poMǧ{�U�}�(9���\Bl9(����p�˓~����em��*�4"�)���)���F:�������f�!�c�Fߕ��]x��9���po[����}�%��@�!3��-���n��j~�]�z)��s��ZG���U��s�u�oSJP�c��P�8�=��zNT�x`M�ȳTnJe~?����y���6�J" =��6�� ��T�DN����T�v�"R�����	�DqX���Ab�)�+B�%P�y�p"Ϫ +��T�yG��>y9�=C���Ѽ=[�AyK�l�L����o��*�#�k�p ц����,�Y����T���M�`��+�M��Y�Z|`B��Ֆ�+��$�!�%��Z�Fic�[���_��L�^�����dK��"3��s��zU�� 3U�b�^Se���hi��G �Q�7SpnIG����0B;x�HO6�+��5�/:/�h	�� �E,���J��\�eu��'x$QM���^�PC�2���@>� CH��e����߱C\sUڣ�/HX'V��ic���\��u7��,�rs<)qj�-*��M�Yn����M�<MqV�2V RU�tb���PA��.�{3�j���
�����N�~�侦���e�X�Y�zĶ���2rɫ�W�^m�D�/��Ǒ�D�cǉY1�ɜY�RLn<}����d��;b����]ª7=��O�͸�A,@GQ�[�_��pʣ�1����`i����'���?"Y�X@ ��0��x��: c��pSa���*��yY*��)˲h����	V���kq�4]��2�u�����|�9��p�Z!kQQOY{RG�΃�n{�=�r~�i�:�a�u���h����o��A5�4�笋��@H"7�6��Ȏ�ۇ8!��3
�r�{�K���uL��գ�U�g˫�O��JB"#��5bkZ�	���o.�.WS�5`����s��աɍ�B0�rܬ���$Xf�s�������]84Eg�σퟘ��e/Ț�7+�p2�����n9�x�4H:ѡ�DM�:bS���3�h8P�}�\�dpҤ����`���jW�˶��1�Y���JT-�X�6���D��"�0D���qR���1S�Rcuk������6��6]U���������A�/���P}�Mo���^�+��ν���NBа��q�3xu��lV�W�@��u����Z���6�a�X��ռ��W�dƎw��ٺ2�V�B"�o��P�����e�</	�إ�ka��-ǧw�� ������p��5	��yC�w}^7=��j�>~(��(�{mEU6U���BE��t"�yI�B��[4)9����PQ�$��'&��?��S!u���W�fK�&u/��L�2�!x5%�ug�n|�o@u���.y�]��)�q2�Bx\���?���H3�2��(2�D<��ݴz1B?��=�	��%�*�&)u�x������>�4���8�+�"���y�i��g� �+)�{��f�k��G����O��0�o[�{�|ucٱ� Қחm�ќ���`|L��o�̥!m/��N �`�1���(�z��H����b�)��%�i����a/�.�_�c��Ŷ8���m��r�L��X�!� ��$;�����b�v	�a�C(eR�Y�N,�b���(���V�9��
��\����ͭ5�A&�"��%��DX� b��˷���-������c�o���F���:�75̇�<�4p#|�S��c�iq�&��o��ݐ_a�	t�J�,��CeZ�.�����<�ɪCMp�0�-�>�w����B?�S@�S=��DO���n���er���W�iX�"��A����M�� �����xd8q�o��#��F�9�
z�-h/�V�i�c��!Lȋ����e��n�Yuه�F���!���*В�W@;�J���.P�v����f�ve�rd��0�����v���1Ȯ��:D(�Ȟ���i��ao���;�ݲK��� =�d=�)}��������=�sK�ƤJc��tSr[Πs�/�k����l�H�Χ��2�aҫ �ޣ�ڠ6Z��X\ӓ��X9Ou�_R�[h�mX/���t=�tnK(���Ɍ���C>{� 1j̺=��ww�痵��ZeYd[�\�?�L:5��ra��&�n���Z�jWh�<
z�'�6x����ޱ�ғ������g�w��o�endr!��E���*����U�����)�>p� H��/�P��l�p�3�8��gny�bZ���_";�r��qʻ����57!�KSI��;-��AaQ�B]M�l�U�Gbr��|��AUp���mݿ)��j�G��Ç۠�
�-�>�I}�.?�^��a�U{ax�^`XQ�9��.4_3M!���_D ']���x������ּ��6�([��7i�ٲ���
�Y�N4y����|����OmL�v37�k��64��d����7_���lɶI�D��|J@�*�(�_��t|�O;�H���gO���D�{��\�%F���nozD T� ȇ�g�ˢ��Zf������њJ���ycS!���{�iZe\�*�k">ðR����	��̩�Ud �5Q�#ՙ���tTф�Cږ*	Z����[u��cW��T��N�IU�����c�*���9	���4�; u���n��Q��|/9Ы�y2w�g�kύ�5�g��?B#!$�� n�Õ�:��?�D>�/Ia��'���H`�KA���4*t1�;�?)�"MPԏ����Q�:�0�s=�wh_U-uޅ�C;�À��g�E�#�Ѫ��7��׌���V��^ �E̾ ���\j���Ǖq �D�X�z#����PdDھ���d+����#$�W�.G�%��t�-'񙗶c�MU&Aӓ��R�X,nh�zȧ�Fe*%�e�l6���X������z7]=��H�*a�a����A4�%�%IL�̻�f.��@����Hi;+��hh����®�m��%M��'Ə��j����~�RC�秄o����#�z�L�	b�4(k^����+i'd����ۣ�t��7�ЩBπpE�|���W���U�AjQ`P��+x�|�Z]�R2k���+]��'�������{8�D� �#s�2�D҅8�<���0d?��yР�Qܢo���6�S���Ǟ���� -+��e�Svx<��sa0*��G��A���w���Ս��)��Pq���V�F�P�M�4��B.prh�*�o�J�8"��q�㈠��q��\����6o;|��X^�n�l�F
�ǆ��e��M ���u�ߓ�x��opʳ�S۞�5���4�3��s(�P=,��k��߭�r����0.r�f�Vx6{u�i�Լ'ԃη4�`���<�9'[יF��["*ȉ�FϷ/�۠>SJ��v�3��6H�m)�|��=4:p�����hSn�q����߳�A�G{�X����j�al�4ߙ����Ͼ��p�4R�5�N��lP�w�M2b_V\	�/J�F��ɞ*�F���B�FB�D�% G�g�VkG������
np��7�3-+UJ5�,���dX������h\���V���x�殜6-$�����JG�'���Xȸ��F�_�	��"����@nB��C&kS��>F��:w-f��9z)�q�p��^Cm[%e�'���3¬g,���!��r��#+x��T@z���$�՗ъH�}u�%�D\�l k㹫��g��,+=zQozR�@���+��Łw���2"94�1?	d����i�0 ������鮊Vm��_�֊]����M�Q��}���w%O��Z+�%!��-H��XL�"�;tv]oz����������'�Q��CJ.!���N���Uu-;m�1�0�.V�S��)�����l�Tb�?�	l�UO|:d�G�n��7�g��lsoM6n��p:7e�Ģ)8Pc*|L�-.���t�K������cl�t��r�ί�t�k{���W7�����mJɫ���y 	}�	b8˓�Ꜣ���x��2b�ƫ��.c�����	�Ҙ�):Q�x���
A�Z�5/��9���>P<+����)a��.[oc�gxൟ��;;�we�ciCs�����R&�$zٸ�1�T2��o�c�!e���/�Q�)~<jg�h������R���~�r����5X�2C�4q�v��o �7��} ]TS��{h�.L(�*��߫��4���K����E�Sm(�Ĉ?�x�@b_b�;��R�a�VCl�*f�/P����r��	�����b2���v4_�C&t���e�D}����оkTj6���-k�wr��U/7M�m�
�g�*��1�p{t�yF�K�C3��!u�x$[$�����x���81K���a$�������'CT6@XunV�Ǖ^�)��� <X�)ڗU!g�ա��<�f���0k�EbpW���}*BU�Z��Fݠ�E^:9�����x�@�*�B%2�5z��W� j��0�m�K�ܻ��~ ��yAV��uuVHCF����V�H�o�6�H$	g����d9���c�L��0'�d�0�Gh��X������is���L�������/�����i�k%�R���W���8���~8];gj%��f�~�!���0�įml�� -�$��|dr<�p��Ol�!� ++@�l��w�ϕ P��l���i�-��;�U�v'�����b��+0�
��KCuMfI�Q��AL�{I!�i�rxPp�ǭP�U{cJ�?(�L�ꈶ�(y����?��H�<bM��n�P��J��-!��v�b�����oUW����̕r�@4? Ti]�S'F���w�ʧ�x�����QfV�ɉ�>�5�6d�)������<�����������L��\#(�h��յ��kV|��6�k�_�1t����1�O�52�9�(p\J�0`UsrTe�@)fT`��]�����"��	�jp�v��ֹٜ�"����= ba�Җ�:���L�P���t��xƄq�*�6J�������۔�t V[zp��<���1Do��3
(0T��Rb��{��T�.�t��D{�+0d�r�e{�z`+���s�GH��Nn��l�F�!���C?]�`���>mz��ȴ��X3�GH*Wx���ƿ �{��Q����0$)��W g
}��E�3s�:~XlI�7�$i}�dH$-���o�S�z��q�4��OrM�ŲQ�6�ۑ �1�|��4��P]9U*^���`�8x ]h!V�����l�5����B9ذ6����z* �G��칧�N�NW�=yY�H"\}5c ��"w�,�kRf阓��!M��;
�������Uj�q��D5�p��Oܭ2u�$��Z�j��C�AD�A������K0��8
��i�[o[���]��f|�r#H���֊��*Oԥ�*��"*D� a,">�B��\y����~�-`�Sa��������RlkEq�X�]�4��;�q*O~Ǔb�n�I�z�4�4"�&70��K�̣+J��e:�,�<��Ck�"r�g�	.{x�En���X�il�1S�Pa
UF�$ܸs�� #��+� Bj�$�ܤ8Q!��Ш������w$���\�[D��о{���:~>~G	�����O���<=�R)���KW�A4���AS��]��^Vl:�v&r�E�B���|�T����c5�)�W�_�0�ĉ_�����E)��G��:n�ު�L����vc���R�	�Lu�ѭr��,���bܕ�ZR-k몎�t"b�L;������p�6�֛�_�Vv�7�Dfט�H�����XU%�)�?�!�1>Ǳx�3W��W���w���܇y���w��sBR���E����D&�q'�����o����mp%r���t,�%&�mx��H]�;��f-�����'��Qt�j�!rҕ�m%�X��m��n
p�g"KҪ졿	�{=��PC�Ύ堦ox%بv��ד,/�(���p[�-!���3Y2S��T]�{�%��;��d��ωE#� ����S�+5�l� N��o������"��������HK"�_�(�t��Ưo�c�<i����)^��]H�K"����H��l�32��|d1]�ŕ���b��??4�����z��S-���m�q����M�.�ܘ�=e�O�E�Ǉ�X��X���cw���@jkI���5�;��Xʆ�-Z6U{����r�}�f��e�]��� ���6	�\�T��i�'�~��c��.�B�����rZ�̽%Iߐ�)��[�(����5=�6�b��4��B{Z�ƽ�鰞f�sSZf��N��Y{��@G]>�ƺQ\Cα[^�w���*P{�tD�C��	�.h¸ZTO���ҳ(�S:xNx-�j����E	�Z��A��6-��@���tP�)z��ou��u��+���p�}X�~��+ƈ;�~gߧ"�,����9	�/���Wp���]3`�f_5P���؍�o�|'�6�D�o�}�(�82gW�m/���P�r�r���tew(�	&�VO��O�8�f$�5�+�����\-u������p~D
k&82��
���vI�zi��)A��þ@ٛd��0��iL��b�&� �}uܰ�6�_n�BJ���\���hu[C��tER�ʶԳ�G��i�9u7�jZW�׋;0�?�r�$/h�~���o���簳��~�#��\6qM��G�GY��,�b¡0���?�_�����^H�ǫkP��b��`ux�V�9=���g�KL��dk/Wr]��`����e`�Cن62�4�y~<�!�;��p{N�C�JrZ��R%�B]�:!��_�iHy9uM��ӠA�	��t>���n�Z���l��c��.�Q0Y#D�l,�ժ��9m#������Dc`ƵR@��*�c3������D�����H0�Ϳ�%�u�S�=�9�2��Z���=r&���e�#��wP���=����:��Ʀ;,�ɓN	+l�����������{��F�_�ƒ�F���c/�G��~�����~��h(I���^�pǅ�����a�����H����lcF,�n�gr��=�I���	��Ueݯ��H��7�?0�	4:�"F��$;�%�
�O�T鵬�sȂ���@����M��пi֋��]���ĩcI���<n�]�5"=�F��E3�#�#�B�he�͂c�^�t=E����!����1x�.V0԰��xd:�����E���Tr����l���f�:�y7�:�aB5v-xz��p`�eJ��K��Q����|N�Z�?��ip�P��N�c���j X������4ÌP���[ˑ�.�)l�T��)X<孚r�B��;�y�[�|�R��(�����5>bBi�,å���v�m�Ut+O�]
Fn�>�gEr���"�YjT�2Ig�PO�����g�t��g.��1ʥ/2�C/J���64��#�pE�e81}�Q#,��_f�eQ:_�F_12?��b���N��@���v�����8�D��̴s�c+�������ѵx�B�2��|��L�~����h�OɌ9-ѩ�r�7�u4x����;�4��p���i:�%w��3f��Z��~���PRw�2M������Z����Y�hŐ)�c~z���i�e���o_�(��1�<gR��ozŨ�Y�.����D�l�:��Cf�Q.�������M�꯴ݼ/�#�c:o��:�$��n}ą���->���'�?ً�����$�*���=��`���%��x�jF�p̉�,����:ʸt	@]b|��m���Nn/F���/���]~Z˸�H�&8B�&�oI��z�[�,+�!�I��*~��v<�R���jw&���k�o;��ZX�V��F`�=�a�9���[6�o�d^c�[h{�潽SӢ����W`X�;l����Ĭ�44Š�h`��0�	K�c�!��=�߲;�I�� mXƅ�^��E�L����3��^bQNε���|YNt �<{U���=}�g�	�4n&	$�>(��Hȹթge��ͤ�x��;�<�����7��f[M{x<gsdc}['�q��8�����Qh]����jn��Ŵ�aK��������' �Ï��Y����E�=zd�QJN���޾ �sE�
�C�>L�l��I��I
�^�;�����t%��:���mc�$5��9�ܼ��4{W��� C��d�Ë�[툉�ԧdxV�Il�"���)�~!���F8�Q��t�R��>�e�}|�t�A/��Y�M������\": ��J�,��z:.~�e9k�?��m��=��^��Hχ���>�#`2V�>Ua\�+zo/o���Ҧئ��o�w���"^<��W��nݮ�_����"X�M�!v�g�|�}k����2q.�u�`�l�2�T��ќ� ����:H}5�� "�Y�V�>����<�M�m��{�E�#K%��l�X�����CH��#�.���R�A1�i�M�o��~�X&�U^�{��X�{���;	��:������[ñ>���}ǏB�Y�G����eOd���;�Nԋ�����*e�!��u���3��+o
[c<��=P���a��ghk�1�plWu 3,�3�t3]��^��RFL�a�~s��H� ����������a�U���nNv-�2?���|�����'�$�N�����T#+ݿ1��%��d��?�!���rv~��u
wǄ�j|����u��	�}3�z9��9��t����m0u.g�]�L�ZT��!DX?���N/w��=M?X� N��%>~��M\R�â��x���0�{dM2�eFz)���?
)RH�n(��P��O��TZB���cD�h�X����ky�E񒷄�~�O	x�X�r��2�g��v����'��3G�^�O���Ĝ5,=�)���E���A;�".�b�n,���P�[�E�U����I��eY\��e����?k2���~����ퟀ����Q]�ɖ�2�^^������~S{�bW]��Ia7\��,Q�}���^g�����3��o��1���U��d�A��7��O�>
���f�w�y/E���V��W �]�#�ؙ�hQ�6z��L����D� �^r=i�h�8�֮L��p^�KZ�@qTv��J������_̟��4}ҽI�i0�Q;,�v�A;�䢲�!W��?vRG�c��o�DN�5��?�CX���p�
�?;�t��-r��1���ol��l2�����e|���n�UU�wMb��b5�ܬe3��1��;bU�M�o���i�"��%�Tiz��~R�ߔ%v����m�5DJwsTy�;��u[��&R�f��{�5~��L�O��t�1fO잋C����^fx�#H����8����V�S�X�ڱ��k�fU+*wxp%�=Js�Ǭ� B�0&���&�ly;NB|)���r+��M���m���յ�S��y��#�ߩPRʠ$�YtJW����S�D�t������+h�u�+q�Vݚ���7 8�@DR]z�8=�Y�Y�9�:�gm�Fc"�L�z"� �*�7.�y��
��.!�K��RF����V��xk��`�%��r��P�׭���*����&׆V�BF�<b�oB�*mW/�"����]=9T=jj{l���
��{1؛�/f�]X�o. ����$sI"��s_�'<��c��5�[��1n�e�7������/�I(�\���(P�Tss�� jz�S���?M����9�q��w$�j9���pz{�3('�{k�+	s���Ӫ|���LO��"�0��ȜP�i%���.�Aϭm�9�:���	ա��_��R3��7�%,�^_���M��'p����5���yϮ��-$ϻL���}�n~oC@5��#)����:N��nC� ���a8�w
}Z��oT:��i��$^P㈮FħIӡ�����-��n�v�?E>��O�+�#:d�fD^m,�F(r#1RWK�ڿ�̡ӌ�(���m��-�ɇ4:�`%~Y�.� )�%0��>&Ȗ���c$lPӔ���}X��n�V����P��t��;"�?�O�W�7FpY�9<[ icn�u����U�,}`�rc�&�m����_S��X��Sm15�<9+���2ҭ��{=��l�D߃%z`��\<��Z��yk��yrGF1��t�1��Ռ_Ƽ��]�(�R
`K1<���A�H[��z��,>�7O �t�u`��Ā{o��W� �|�x22�����(=���H��-�e�P%���/��4���̕qj�8)��u3:��=|Կ
�knk����O�ec�Q�BM=gYTp��j�Zf٠�Ҟ�(�i�s�~�FD<��V�*�G�21��PT�ja���p*l8�ݳY��18��ۼ�F|}�PVv]���������Z����D�T%���Ӌ���)]��WI����e6����ۻ+����2�{i�A��������]�m� ú���x<QO�]��7C>�GKwh~���SDjR�\6欽H���M�  ��6���cM�G�P�X!A�(i�[^Ú��x:k�Muxy7��� o��:l,LLR+3j�]C�[���Q$�`7HTȜ�X�S�<I��#z�PDo`�:�:��Jr��Y�$�����ʱ����A�B����Ct�L�
�eSW�#��ԛv��S����px�m?;;�7-��o6��㢱�I1��hbn�NW!��m�D=�[%
��B�+�?4g[(y�N���R����Oev�>�J�������潭��|������'{k���P�u�}4m@�Q�]X�v�QB����1�%�r��t��������y]�q3_1����=����X���U�Im+����vT8��w&}�Q��e�G��e��mn���umt��b3@������@�&���)��L�
Rh Z�.�ߛ�����]�у���*@JH�Y���X���}2V�Ƅ�w*(�aN}�s����qlo�u������y"}/,s��#��M��V#�gZ*b��"C�랠n���_N�f:�M�?����"���irqUku"/�ha7��R��Ԋ�$��m6K(�A�<X��;4;�a��t��^�k����UҞ\j�p��~��LƖ�i�R�[6c+�������u�#�3����
� ��T�ͱkJ����	��%f̼����_'����mU�6�MciÙ��,�x�DG��H�~7 �+"�������k+�ډ-�@����Y��`�S9z�sǕO��v4��b"l�:-,4�:��4��*/��YK-y[xUAc������Pj�"/F��ԓ���J�=���Sd{��))�1�b��a�E�1����a�Oa�3���P��O�I�2�5PV��B�͓s�s"���4��xm�~`�T����2��gM"��lhXV�[伻���ө��Bo��Q!��5ZP�% G��������ʢ�2����d���>je���;[�OO�E/B<i��(H���7w�*߂t�`{}XFp@e�o$��]*�2���Ȩ'�c�E�i�l�,@	�i��dS�>��	�+R�����
	aI��>��#��<*E�oCJ* �6���Q��[�wF��y]	��:w-�zUi;rd�0���*S�EmT���`2e,xW$H�� Rg��� #ڀ�`�[�Pw�nlن���<m�r�(0�i���(��R	�.��M�rk�C��=iʶ�
�f�W7�Ί�|s�6c�W3�?�0�}�|h��`����ŗ�JTt�婐U� Qf��xzH��6��>����~q��. i8�e`��ν,���0~��[Ȉ����/\�ΣK�6$;Cr�%\p	�i��ͅO�MRX�]�p�|�^��ʏ�"�	��kM��	I�T�!N�"=9��S^��f�=�
�QO�0�%W���D�.A��z�>�>d��0~"wί+K!�u����b�C��lz���b��*�ꅷQK�j��}�	��?>Q*e%���`���2l����؆���F6�xѦ�Hf���)��ʴm
X��m#�hyX�Y�B:Q6��A�7t���G�ni.�h~�=1Mͩ���Z�=q�w���LnaL���[��$b[�H#~1���Gb���r�iR\#I��a��R��-����;Y�|�)�sy'�EODi���-#:��`��dp�{/���	i�m�:�����g�ӫ�L6����Uc{�(n��NDT&����f�����i8�� �')>;�7�hU�������&w넅^1����~��4��И]�g�\��^ ��/�7��{�S]���R�g�>&S4��dm;�>H	�V� #�N���U����J.��A���,��)}��R�#L��Jt�{�r�$��		g�=N�n��\�.mw���My
dDT������Tb�A�i&����y�=���8��\e�3[�ZcM��~���ۮ,0�|�z͇{Be�z�{�~{x��:��#a,J�}�\��'��?<_���yU߼7.~R�|Z����Aéqt�Y�����GE�Tm�jw*�z���g,~�t�a��Ӡ��}*s���.Y�Ln�b�ͻ./X����	�nF��q�4���d���hv��OC�����U�s���bnZ�iS���˩E��Dȸl������ ؗa��Wvir�m�0�3�Q���~cf�mv��E��)��`2$C �˳�ܻ�kRB��wF������~�7��C�1�| ����pT�j��ɓ�tӳ�m��
�w0ԭ��S8ט���M��r�}��Ÿ>5����va�yj�e�������F{�t#���"�bt�v�Tl�49�fWh��h��R�*l��C��y��o��瞣Ϧ]��ڍ��^�6�X���k���0a�����ҍ^��X̷eHb Q ��$A�{�F�m��aGn�vF]�=�Y*��mh(OZ��3���v���	���>�4
s�q��5�5jf�n��k2�O�Jwe�1ĸ�R�O���:q���z׊ĠH'�.�E���)R �P#�C/K�8}�g�Bn��]�|ʆx�G��&q���>嚌��"��'x��QT���편��Nz�\�4+�B�W
2ac"&���8���x?��,o��z���O5����2%��H-�n�R�\�b8� d�z�C��8ͫh ;��g5�
G�w���q������XS4�&v���r ɚ����K�<U{�Խ��{�Y�P�E�b�R+SְI��s���Y3
AS�u]7�W�xԂ����!2��e�-"�[���wg��m7��{:?c@Ѓ鮡d���\�9\� 
�nz�5+��\��#@���;�s�Q	���!�h��1Y��v\��8�����Q��m�2�ٻ�H�6ҹ��)��b�ˬ�,K*�P�鋒��W�	p}r�E,ǫ�E|�[t�����F�����>� Z@�x��G���qLܲ�GX���A\������{R�-�����ֺy�w'����CQul�'T҂�a���`�؉N��۝���~�i��]5�3PB��[M$5�Ϭu%~�!�p5�!F�Jz�����v��ˊ�ǤK8����TMk���EL��N��TWs4Ո�7kc<��{!s�+�l>A���?LM�e�����R����ЌX��~��知{%�P�q�N��3*R3�%bF�1�cu"�%W���-*�.�W-�U����IR=�J�=@g����v��C�w�ܖ(~Մ��O\�w�l��7I�����M�n�� �y��u~b �̸mv�(�ox�߀qvnJ�����xp�R���TLR y�y�M�pP��[ �%��Pn����}y�"�$������:�W��A��[���`�e��܉5��h�H(`mQ&���c94�wbwy���[R߁G֮���Z�y�y޿$��T�x}� ��y�L5�g˗��x@J��ۻ��/.K�k2n��H�P���a -M�_ܿg��z�����OR�*vX�7#��t�-X.� ,<�t��b�;��R�����7�����t���8Z�ńE�oHP�MJ�m�����o�تf�Eސ���#;�'�Y�~�{��4�������!%ӧ=�ֶ����N����-K������?;��B��T�7 6�t,o]�Lb��^M/��l��a���.n��M�����F��C�Fزn�vY�e�{oX��zZ����N�c��tnY��8y��v�걌z�Q@4�N�hm�9H	"�*Pm�n��:��L�(��hr@51�K|ܸ�V���,5�SNt��|���������z���>��`���~=QH&�I[�e8��Y���sHQG1��8WP����e2E3p\C�E�ӓf��������N��֖I_��@�,��%��@p��(E��q�E�}H�v��:@Tώ6�9'JD���`���Il4��ؐ��� g�X�>��F��.�����5��=���sQ�v��	�h�����e��(ǂ��
:�9T���(  �����\�Վ��Q��B">�U�3i�Y]�W�xo=�J�5�}�[��?wIςr⚕a��o᪻��Z4�����8�$�q0=�Hg�Y��z�jnZ�~s̹aa��j��&(�W�j��ή�	MԶ�,�Ӆ��G�E�Ϭ�$�ԡ�f�,<�����PHR�ؿU� y' ��M ޾(V��Ce'ˊNK�%������A{���ɳ���B��C�i�!l~����r�뱘�39�_��P�0����m$����C��_*�Ѵ�{
 &#]�6�N��`�]7>����V#y���ʆ�c:[�z�ԟu8��.�b@G2e^�J�W2��Vn��t�S}�轍�b5ɿ����N��~�j�X�<�/ʜ #
�aT;�٥���Y��X>nSq�66(C�04����ɭq:������� "L��<I1x���M�CnX�rq��Mv�En?��~i~�d!�T���]w�$�f���� F�3��zEOf���XyPr#(r�G� l����Ho=`#G��Ѷ��O��ߟv!Xb>�8��1c촳�LmQ�8CML;ůu{�D���t�H*\���{�>/��9 �9,&2��
9ÓB� ~Ƭ��;���PUd) �`@����h�HAȡ�[h� I��A5����ß�/0j���YnWSK�Z�U}�Rc��ھ���x��@��/
��;Їm�~��/��X�E�������G
n�M6ēĝJs��ƾ���ʜ;&d�x����M��J[��r `;�֒�0WZ��H��ɀ�k��o���� ^�^���]�����ŕTY;��
�z-�I�Ч'ҡ����߂vZ}��!whI�Z�_�8;�)�%gv{�H����TK5�E>!忿F�9l��
��0�����Y9�&���׼	�����r�}m��g����W��G�Z�W�t�\������������e�K�vS���K�����f�F��7�������ȣy������\���N���=(*RZ��9]3�'Nh�	I^^�@�#_~�g��G=��ⶴ����'5g�z���Ш�H-3����i��q��j��b�!�[Fd��5)��kđa?�C��*����`�M7X��2��W`(�bDXJq�Ǻ�g�l���C��=RjPT��D��~�~���]u]���r����c~+�V�,�r�06E-Y����XCU���M�s�n�&ͤ4�����cB���Ő�>�C��#L���E;G��M����#.�����%��2��/J�ϭ���&j$��*�|����E�+�1����:���(�����J�m�H���
ކA������ P0�^A�g9_.1�g�����/�f����zec���:R�b�Uud�)��&��el�8�cV���;6��pfO�"kW�����R�c�{�t���ثen�8�IFO֪���lm��%�9Ma�$9���Ɗ�Ld~��k��/�s#�xe��yP���z������/f%���֗<Ƿ�:��blo�����hGA��f}����#'�"�m�F�O��F�k��ES�T_mi*}H�4ey(�Fxb�<摞�o��+���C��L!�9&��Ũ�Hl�ǲ��AZ���dq�:R�\����S�ϸ�i�ê���Σ��v�eÕ`!����ī�%����܁���K���-���D�o�1��T'7�-y/���q��ɬg꯵R�Vd�B�qXaj��JӠ/���"IU�xsl�E��	�Qcsǚj�U���)�R��etL���E�1�Pĳ����"M��ڛU��ٶ�mM��Ln���V�U7'lg��b�%W�����7,�?E�9� 
�\�Jɒ�]5w�x�Z+6)T��l��8󗗛�4X�!����x[��/W�  U�g��歴Á7��G~Ƈ0� ��F�3ט�4�2I���zAr���C�3������;{
u�t!>Q�d����_Ô��23}�tpH2Y b���Pc�d��dh�S3T���@� �d���&���0��D���~�s��A���G@q�J+N[�?��	��k�`8s�Z��qB���5qX�����LG�8��՛��(��E���!5���h�X+�JB����O��Y�Åw�˗Z��:i=QMQ�:�4[�(nC%���h�����]X�_2�Q�u����&7�Դ�Ɵ����ZrNL��i�˃v��QD��2�;7 O�6�E��F��]zKF-O�(㬹�3+&�9�"i�F�}b��!�	D=����g�[�잃_	��bN$5D;�ޖ��iV�~}z���9TNŸ'�D�M�X�F��I���E���ݧ+� G����I��t+�ѥ����<�/`٪�T}#iRٓ��8W}�� �9�e{���k�p�l&"�a�`UI�;//�ڻ��8����f��o�HP7�Ʃ�t�)�YP��U��[�G�v>�C���&�\��|㟠^Mכ�����j�J0���t{�m�mIP,��� ���h�Dv��:��2�?�[T[�Y�W�&��U&3�I�Nǋ
w���`�مD������vJ$�/��p9ɕC��z�O�缰,�ע[6 �s��gE#�?�:����C�>[����_���ȝM*���#l�A�̳�me;6�PͿ=��Y T|*����L�� t�lо2Ŷ���E��D��l'��~My���
�h����u+h��#�b#�&��o/�Z�z�Ì-�L>LN�����0�ʭ"�0{�)�n�Uue��S�WA=90cH4и���-�]؃�1��7��r55dr�q����"��i�Z*��n�+*6�[�8T6���
�I�s֟���m2���*$g��U���J`��)���W@Y�2W���<��Suk4*�m�l/f4L���ǝ�N���ɣ-V���G��.�m[\����<8X��Wl928�	�jG��R��7��s����O�1�"?��\����  @��������S�gD�:P<L���>��q�ݓ��YZԘ�[] ^T;�<e��8/8x�5��,�M��`�0�Ɩ)A���3��j����=�+��R�,�t�w��щEu�4�L6��i[s3��u��3;#���^������b\�e��gw�_K������&'��U���J��[g�맒7��%$RP���n���:z�����ku�W�h�_]l�"�A�.��;�9�Es_=oX�c֩������,p��/��~��[�y�xc���夼`A���2gʃʃ�9,e��q��Mn�=��c{�x@���^|I>n_s��h�&�xPQ���CW�Z|(��������sʢ ����m�ܨficᏘʔ�~��X�������%����i%R��q]oE�A! Q�L�����@���Sfo"���
����Ұb��Kx�C��Pé�v�s�(�<F����6�J��zDBF+���خu���Dи�â����EJ��W1
�'#��Dpc�o#��|����z52ȧ��d�,���At*����:3F�Eeh傰G7r32�[�G\�AqWU��9g�\\�8N\[(�)��a�Z���.�]u%w6l�6d[8���K�ZE��>���D$T� '�⠎������V�Y���zh<z�ĉ�4�.�1fM�\㽥ɮ~���C!�{kH+����FA�b[Jס���������xf�'�7*��n��7^�F�V[��bp������ؠ�`�=��~�ң%��H~�>�p61��F�0n������=��� k�b;�DJN�ap���2�j��2�vjV�����jԦ��s���G�{�).5����!r$H޴-�qj��m�/D�o����?���Mf��؇i�a�n�ҥA.��e�L<����2�^��O�t���o� y��pˇ���[L!��A&ܧ[��S�:4qo�L��$��ֵ�d�Bx���dd*F-��IoT�𭈜�È,6�V�~���E� �D2�E��S�S��f��2����	�0z)�� j=�!��Ǐt0N�fs�~���� �3�)���
���"��Kz6�T���?���^6!��
�u��j8�v�v:}�­���l�!t�j�XT �w��~���l�Se�� �aȃǬ�<_f����c����_̦�T�LL�Nɑ������G��<
�����S�_^�[`��`�Հ?����"I���*���L &�s�Ϳcz�r�S*l5�x_�/�}�X��fp/�M��(�ޒ�9�I�+c�C���%���m��#~Q��9άm[�����M��{|`�9�*����+��>��j���1�����	v�A��Hk׷��rn���f@L���~�qɲ� ��U��c�����G��M�1��G����~����ǧq�i'2z�XK��+����ݘ5	q�j˛�n5L��f�����V�	���V�zc����,"�Ky����<a>
 �{[��>0�V3L��ոOH`�iӝ<%�N�l5�'PGbL+�y� ����LfU�jP�ڳ7iI�~��׷���= ��W>�x���u>�j�u��(7I!�U����ٗ���(�����(٪�r�,���'K��xGi�}�(����%5�{B�q7S�:��J1ZW��4���؊��k@�º��ۑ79*`96&\ꌛݒ��L�93�8�-N��0�D�{�@��]���"���ʓ��G��t=p�ON�ɻ3���^N��UŰT�y��Ŗ��Ё���I� H�=�H]	~����w����ۚ�^�%�ۤ����<��d
y��&QGlK�!�ƹ�8��'� ����FrOj�݇�H��?�d��Ffp�3���*K����o��� 2M���+� 	`��U{F���L�H������n~>���^�6k�;�{;!��/g�����7|��,�q���ys�W
���@Ð���i�<&U�+D��;�A�2�!�,�B��Uf�i��jS6�;R~�}�vn�W[ךF�鳎������/C�DX2�������]��W��B�=�h�P�]����٫}S^��ay>��~���ը����9(ڄ�FO�u���3��N��}f�����I�x8+���h���J���u���������4YZG)�*|q*ó7����䬉__�O��8d,c���I�]f!I����@�_�}��V�}0_~�n�u ��coU���z��	�P���ؔ%�N��Z`���v��<�Pf.���1"���oU�#n�殥��?��;�@��"�;�ñ�#�2[ڢ��ވ5���W����fuy`�?]p������]��� t��1&f���%���t:��B����8V���,���O�϶!�q�����NW�AO�;+#Yg��.Xgxi gdWr��@)���L�
���6�[~oiV��Ż��Ӡ���l"R���Xq���I,ď
\t��l�"<þc�n���s�c�E����y�u����Ǹs��a;1����z��im�����|ы� 	�U2��ݘ��)����Z�x+���E/�.���Ѭ�!b��
Lp'T�_������[���	��0�ќ��<T7>��g�Bȣ:�w��e��v*�X�`d-V�Wn�R�#�q6���_�A��zOy�*��+Q}���
�!�7�Mϵo~褘�!�9:j:�d����Я+`0�ݟ��|�®A�,����ѣV�¸�Q]��`�*-�D�Oȁ[#e-Q-U�")�3�P��%�}W,���,nd)�r{W��C�6Z*@d���B�������#��H�^c4�ᔻ]k���dN!�R�X�	����Ո�M%�j����܆��D̞�TU��el�(���=�s��H���*�����pQ�x+������x�ٗn�}d�&T�[�O���X�a�ڪ01��yCc�{/���O��Y��o��*p�o��P�Ď�Pw�'f�?�t�x�����q�W���A;�H|O���Je������%t�STd�6��9j^c�iF86m�ӣJK�y�M�e{�:�r^��#��E>��%T���?��^�.���X�A떻���m���������NL���k���t"��W�T��S��h��� %�8��̾�h>I�])7�x��A�H�tR��i���i �ZO%Nrr�������TFMh)�r�b)�{�"���C��Ǽ>�����*� ��#E���w�ޙ9T��ST���)M�*��ku�V���%��w��{Λ�e�,� ���v�M&y��sU�"yǐ 1�iy��6F@ �f5K>Bc�x�s$bX�)h���]�Ş�%�*�(���-K�S^�I��Q���k�1K�  �|����[G��$J�
G�J`��Cw���,���x?Q}@�qr�uP*	�{�RN�u�K�X`I��m�Qsn�n �ד̭1����Ƶ���K�/����_�E��2�狦�w'�%V>
��Z�� �Gq�	���C>U����_���t���lSq����P�+1�	m�,0����i��c�̟j�P�gJ|�ށ�&�WXO �&���mO�N��.%�Ft�>���`oW�,@2tE<�k)r6]����40K�~!P&�
吪�P��|9��b~���	\t�m������aG^�<g���hhൖSӯv/�:�AmCb��a��J|�/��R@��R�e����A �d����
r�)�b^9��g*X3��6iI
l��5�P �o��d�����uH`M�?�(�u}�T���:����������Y8u�v? q��f�����?Sfr��:胔U�oxǆAy~��ԯ<����Ź{�+�>������[2���[�!�#�[�͕ X���N�e���W6����IKy�V�Ғ	�e�9]�z�Ū�p���}�%�/q����>W�'L_>���9�f�>K�͂�1⎵5,��O�s�����h��N~��Vy��I+"� %���g���H�˅�xu>.�bKE ��X���plU��W��ھh��޳��Uh��=���<�Ac�'6�\G�͌,0&c���|F�i�9*H�1k��
cA�٠�Ydc��	b�8����� ���G���Ŝ#�����X��ma	�t؄!H���G���b�I��i���{�+.���;��1����g��[sW���F����
�x��˸H�>�
�ag��g�ܰ����Qu����gS73 ���`�pWW��#�1A��[�ʾ.5�t�m� �<%|�sq����V5ʏg�*XîJ�q�/W����֙��#�K��MZ�?���o��_�J��蛣bH@�'TK��?S�	�I**��o�c}�������ܒsU�'~�們m�v�]�|�6]�^H�����/��<7���/>��Q|+r`	8�,����j!�ϣ�Z�P�Ȟ��y�9�MT3����%B��&�v�sַ�.�l�&����gؠ��:��1
I���N����º������6cKw����¡��#�k3i��I�óA��i⠗%)%�Ω�亲@'�>�8X�|����� k����6R�([�?�5��(&lW�-�X�J�o@B�l�Á��϶D��׈������"ou��mn�m�u��'���"4���D@��c�\�w�m� Q��u�[A��m��׫<�`VQ������^LU���`����;��=
f��OәI鶸�UY���<�$G;t�V.��(v��cʁ˔Fs<�h��G�*��>��v��Qj���L<��4�����q䋹[���2E���2�72_J	I��F������E���$����'3cD��$g{�4QL;�g����IE����D�y2Դ�S�q�Љn�X���0��,GEŠi4�A-_+Y����Z!���}�Iނ5"��.�ړ'о��_Op{��%.+��/�i�y�,?�2�'��v m���{����d�Ð}��ޣq|�k7���~Ot9Z�i��}�5�'��^1KޥL�8Ço���VO�� �5�6p�#����_Ե�^��ӹ�U$Y�� ���$c@a0A�Q�o�Î�Q�,6��/5�r����}��Gg�e�V^�,�"��)O��(Jq�d�)����p��A
I�*����|T�Xnm��OԻ��Q>���3;,O�隽�sT�"R˴�L��s�F�II�����4���BfW��ݢ���P�%M`�����q�S��),`bra � �:W�&)F���7�L�2`�y$�q���Ȃn�z�{��C	N���6~TC�����ƫ��$󷈛q�u�iˎ@:U���>�������������B�vH²�[3cJ�
��8(�d'�����*RG�C�����A}����s�	���bj�f���5^+n��V�	��C�e�w��a��\����S��v��^�Q�-�[��C���v�VB��b��
�$%��������k:Pz�+�,��z^����;:��v�4�񄎄�쯴�ņtu�i��L�'Ԓ�� !�hE�R;/���"�𑋖�=	�\���_�Q?@U�抵�? ��wR��Q
��'.F����ʑ=���;�Aǎ��VG*�o�ޟ=�I��z����R�U̕��R�Ę7	���U�0|��{
e�5�v8V~� �t��7`^���/L��.� 1��r�T^N��0g�TfH���z2l([�S��aZ���H21��Vs�@��bw����#?��ڼR��lllV!�e8���\�"�J��o��l�-��k�6��R.�Ɵ��o��$��3��-ӛ��h��hJ�.g����_��VS�!��A�14�KU�p�/EX撿�jI�/�YvEb�D��<�r������h��W���\�HY<�]�7��e��v9��f˺}x%{x %UzH:�\l�֭ߟ�f*[��&U�o�g�Zԁ;�Q0��S5���k��+m�W�7@9���{�K7��{��>2��3����Nl���7Sm��v?�r�\�oBH��oJ���f�n�d�&ec�V�,z��'.���et��u$5�s �8I�K�0����U���oF�~6�d���25� �G;N�X�^뎪��q?�0���=CP.S!��I��H�"�d����Dg�{��+��_���ꌂOU��l��B_�$���l����?��-}����)��h�Ƥ�f�w��s�T��*�
��j�O��^_)`6���i�;��t����%6%�w�V
� ����ʮ�$Z�9�C���e����T����y��;�ġ��ҧ�9õ)�;@Q2s�	��D^�BO/`����[	Ό]4`�x�J�_f9�R�/wu-Q�-:�
ٞ�I�N����&нU���� 
�@_�aS.�������XPT�yv�͹9��N��zY��#Z�s kO����c��i��HM6�[��QPz� ���^{aE�pWZ�����u�kn�_�)5|j�91��+��!o;�ש60�^+y����9�Rΐ����^�����������Fa��=�G,i�@�\��3�H���#�s��B�u�/���m��>�ݸ�%IG���-�xg$��M���paN�� �9QCފ�ķ�<����C�ȕc���:˔aQ�,V�>�O�8\I�!7��!�� ����эz@�;�jO�)8Mw�e�`
�y���.㣓��(�{�c�����Z�1�p��LVA��ҵ&~JOM�BJ�f�YZP��x�$���j^�h��n΅E+Iq���6Dx�q�N�Ʀ��a��_/[s��o��!Cchg������s)G�ߝ/�!��d������ύh��a�Ȝ��o�Λ��~��D���Sp���cgi����^{xr.I��@W��9 �E�кB7k�{i.+(DV$\�=-2�R�,Z�}|(R���D�	�)A�[0[�3%	��b�{ֽ!�R�����`�9?l�up�O��|� z�m�^5�z#�ǥ�ك5oSpV��v�H��2wC�+����$8K�E ��[X��6����L���wQ�D�稐�WDL�q�}�gd�����<���z�)�]�*6\�zׁFL#w��+�e;�^($��^*�R8���LE�WŤ7T+��"��fK5|5�T�=�!Xe��#����C��7IZv`�r�|6��o��>Z:�.���g�v�g^| �"�FM�. ����gK�N�b�R:��(}�h���$�맦s������Ϗ�#�2z�|u;x���Bu	�*2\Ⱥ he�j^�C�5�`��Jk��	@63��:��)+�%�#��Éf�|�w��<+�&�6P���5�d~�`$��y'7�؇1�V���` �K\�Rd��:��[���a��~�	H;Ҭ��/x�|/�:,��-Hѕ�hۜj~�nz�jF.���|�ҽ��å�o�����%87lC��+����-�`�fW6�������q[R��H����o�):���u�`fԒ!]�W��(ق�cA�,����>uU���c�|W�`y�U��v���*ǆ�\�k� p���7�WF)�j�,��(�(@�^E��=�o�U}�b:N���|�6Gg�9NE(:+Ut��xFYm4t;�8I�	�.A�,�@�u���`N�@v5-��`*��o�ibW6�.k��L3�d��u�Pv��7�{�EL���F�J��ܶ�ZN���b�������H�ә}�!d�~V�=�v2�C��^���(���3<��Ȓ}�uI�v�Y����bi�O��Y�r�؉�6�PŧaE��\��,���sac��~q,\Íc�g�hp�j@��&��&�&7&��d�r��PV�jY\j�H��tm��Z��� �"�=ݯ���Oe%�!^R�=Y�mqΞt;Z�T�AYǐ�|v�i�����#�`���pg<�b��uq|F~r1�����JI��V��'u�w�Ԁ4_��2��P6�:
�C3\	(��C�5z跩WQ��g��j�d����}`�}��sD>a�:yR���f�c��n���?��|����+�N�$��&D%*��̪i^ݫ%��`�\��{����OjI��A�ɆMN����U�z� �n�0���% VT����ע�}/��PpbDD�a��o���)g��v0���mB��Δ��ޕ ��]ɐP��� �`"�_]:�F 0����g�\�Ci*�o���'%=KI�ϱ��� ����G�$?���H�`�k�2��DiY���Һ��i��q��m� `�
G�bpH-i�?���{fnI'Ģ��OR�wc���u%�"牊������ �7By����}��wn�!��ʜ�S��+������	������OU��(��Z�-���]�5� ���� ����~uG�.��1�ĺ��֭{~�x�'��>X���^4�L	�F�9� ��}t�d�C�K���X��Q�	P�J���B�E�_��T5��V{��a�^-�p��+`w�V�I�Sh#`T�B�~�+E_-�t��*:.P����x?�A�A7x�z��1M��Z��	0�v�5�ӉF�����lyx8��#�<Y��Z�hPW݁)m��-H&��њ*����`�4b#*PM���$�u(�r�(����6�@�WSRY��U� �|a�أ�Lw/�}����,m�Bs�?�, �7��R�/��_T�r�,G�tA�\��6\��C����sm�D�\n���[�Bc.�s��<m�Ǻ�Һh��)S��������뱒p˨vs�x�S6�z���]���<�ya�.x�S��6#�+j�4�3��r�BY� � g*K`ב�<>r���m�4��0���|�#z�m�����Bᨃd'��""<�r��zө�'�j��䴠�Ҕ �ݸ����5@��ēA6=�bz��a�N����s�A�y7*��r���o��-����?�!��c�;3gY<@�M<���j�T�4��?���Y\� }��I�&��qNu�b�c�4M��T�m[v)C	���u�oF��o7��X�K0�V�q�����e�#Q�a���)��J!���ƜHl>�R���V�V��������P�^Ջ�a ��-��\&e���&��K��ȴGS>2�x��[��|A�� !L-�XW����o��b#��-�1�����3���*v_���F��Y$�e(�[��n�d$��k���1����,B<K���#T:UT�7�BX�>*�2�)������؊�,�=B�a�:TɣF�)S�b�@]s�9��`�c�c�MJ%⥇6�)�<o�z�vЧ	�J�b������y3Y �t�5�����c��S�#eH��x��ܜ��WT��R��!6�\\E	�@��٨x5+�Ҁ�z'q�� ��B����O���0��T^�ⱟ9\��6�� Xr��['6����Hm��Yb�{B��TG{�H�Q�]W'��e^劻L�^RP�R��iY3&��
i���$z�7+TK���p]۹��4ː�_h��� GsJd� �7�Kˊ2��H:�U�!���t��G�7�P��gQb�T�֏Dǉ���7�����\]���j�~�[V�!�Y��$��-�D��<d��֭?�Y�@���~*zJ61%��K�\�eWӛ��h����J��
�;뙜#O�" y�v��(�FS8�8V2��Fd��a�.�2)�G�&�8Q���\�eˢk%�8k9I9T6e���C>y�dWsaA&S���ej\��E�ۀ�̞Q]�Xr���z7u($�ؚ������Җ>�W����OMn8���쉲��3sn��֓����Ӷ���	&�����#A��5�K���DyqlG�|���A�T ���s�6���ܘ�okE�B�!��f�R��L���Z|��M���LR��~�����4�4iJ,k��Z�OW���ŧj�EٶX�8Bw���4����� s���ȦY�wK}͈>���!Z�_�<A�R��u�K�D� ��h��b��}��o��'(º Obo	{^��c9Z":��!��z;QK��=S>@nH5���_K��^Q�]��B�h�5��jz�ڻ
�H7S������Kfl��:�X�!��w�&��a<����wF�&�|zl}n�Ƨu9�\9���Lu-��-��ac�g����HT
E�j�O�J���d�T.���x�Ձ0w��W��-��s��\J������ھl�9ޕUY�����3��./m��ف#Λ��ڨ-��Q�X�W�������~�A��M����a��sG I��)'N�v&��x���6`ݟ&#�TCxX�A^�WA��c^�vyu��؞r�'+'����]�h�eN�b�q^���}��I(!5�����Y���Ѧ���ӻ��o�qC�y&n7osaD.̩`��D(!����6�)����q���y0`
��rP�YQ��TZ�	I;���?`�%��S��[�Xa��4\�×"ƨA�x�p���$�|Ge4�2���k�'֣�۰�x	(�9�IwC ��rn%|ƾ#�H���j�S�6#�ꨭn
���F�|�� =�黤��7OPA�1�O�&�#���>נ��22�V�V����Q����}�,�mRn�kxegi�m�����8'"�"�����׸����k��vcL�g���>��;�6����~�8e�ԸT9"��m:�i+�--�2%,�D�~�h��"y����#k��fU%fƪ�G�{�-�~Ձ�������6$������,�D�J$Q��������*ܬ����w�`�������E���\��uZJ��,@��#��x񜄾�աf6
�Rp�ا��A���V��Q�Z|�/Ka����A�j&��R�U�b���3�٠[Ξ����[L�Y0$��������_�:�s�>@ {���I�����(ݞ[9��7��`�U<9E���,[-��.�_}~zj��	����ߵ.>��\�����X{��ή�I�
�LG@H/�e�S����Ű��/9~�qj
���p�R��9�M�����:���i�t�AG�a_9� P����4�'ܢI�tؘ2ʋ�2��AUn4� �e�&�iҽ��j���C��y�.ā#�O~���%��?�O�|��6|F6V/�y����	N���_�}�o����	�2G���9,��^W���CcT}ǃXZi�?6��h�<y���|��M�P.b�T��=vM]y#���[թ�"�~Fi?��r(2yU%�Z&�/� u�3�8���= �t�iηp�2�n��������0�4v��<tz�����	^��u8��7A۰ad��cś��u�s���dv�t���l�Y�L2��n��%O55��q��#�Vj�:�m�11�ꑆSkl�8�7��<����r?���X�,�ID�:>���'�-���l~iZ�:���8S�
�[O���k�2%#�V/�\���LEc�� O��7Z�<��ʙ�|�q��#��Ȅ�P�-�f�;�d�H�G&-u6�C���P�1ӝ���%yH1Xi� �9fr�4�(��`
��h��>����O`��)�W����7��VQhAo�����zB޽���Up�%���ѹ~�W�Ԧ^�m��8h���e�|�d��6%u�t4�>��j�Rs_��b&�'�X�Tf2���Z�#�zz�B��'�x��_}�0F��U��WA���������X��	n$��)M���a�T�|��sYmB��B�����IF��w����e��l��8��X( QQ�˕��<�j�J���� �Mꋍ �>���h�	U�R<���pp��y�kj��i��輑���ڽj�f2 �~��dx
$f������n���b䴻���8Ki�+�U<�=W�=���[�x8E�:�a��܊��+x<*�W����n�O��K4a���I/��i{BmX�k��b N;�_=�]	�P����l����y_�X�+@Tj�Q:6�p[X�ޮ�Q<����^%<B�X�l��) �U�Oq�����������'S��N,IX�	�<�tH\5���#�����q��EV}1ī`�&�IJ =#���ҁ�v�Z�NL�P`�
��Y�d{�i/9�A��L.�{3ة�ON0����60��h=����RX��퍝�(�5>��ݘ�F���A:��Y��g@j鞆�bc[���<���<��z/a~�u(��}	���w�[O�:e�g�ǆE�s�׽{Ad��1�S�����S���
Lr.s%�z1�5j�ipd}�&�ͳVO�V�a:/̙�a�����o�.�8_���km����6�Ɍ�@3>D�i�Ě��Ta49qoc�3@�[��C�ts.�ȧC2|<����̍�E���ȕ��J�ХQ����4M�w�/�xY����N6< ��è��LW���]W��y|EZ{��><�f�K�_
���d�w���V���g��JNr>�qI�?����nQ�l8���Ú�?[���R5�����t>��
���f�<�.J�-�r�fd�K�$��Sz���}��d� �=m� W�d]�Yì���5�;I��:+����`��<�jFo�ۏ�l�����
���<EU�¼���DD�(m��y=�)�`ԏ��a����zByD�������8Щ&�`TAXoT���7?p��d1�)|��j�D�H�������gfjC� ��H�M�DW�&D��=Nʼ�����I�R������rz�6�6`s&b��XX�\�u�7���\m
ö��P{�h�[�ؗ�zULD^l��/[de���R��2���5��h��޼�΋vͺ~�{W��v��o��jڐ`�oCj%�rE(�|�v/�3�8*�8quG�[�tX�߾�dP&�@gMќ)��ά��>�v����� ���4�������\%` @ ���k^X*���s�/��4�N�c ��H9Zb������o�4T��r�@[y�\���+�����a����^��ճ��t(���^��x�TB�T�ҍf��XJ�֚�g"cL�2
�"�Z�O��s�R���wY����Q��^I��顑'���BQ���
Θ���`ʻ�͈MN��U~��3#,��7,pȢ���b��|��qt8#�����+�sߴ�-C*�.̐�����)8��Z��Z�koN��/5�eg�e�9u��'T�k��E�p}CHL]pf� �(��s>R퍕e�B[!{D�����N�><
�>*Ua��j�=>��`�,%�/�4�ޛ�	��S��o��Տ!���S�>����s�5���
� a�/\(���`o�/��{����c1�ǿ��O;{p�S8�J�k���.F��bNlV堈V��l-��A2�4o1��@TdӧO�@�n�u���r��Z2ʆ��̖M����`��m��mLCa.��s�H1jC��[�J�j>Z��*�$�?{� �r�Ҡ�Ӵ�1�y�s���n��3�m��u��B��o�O��C�eӎ�n�1��:Ʃ
ӈ��wG��V�B�$Z�z��n�m����2���k����5�	E)�r�Rܒ{�����i���?�x'���r��K8\���S��)a���^�;ɻ[Su�̩�A��a�M�߷�/�/\�������[���6��q�[ۻ�9��
<08~�*���.A��&h��R�ۆ�&nѦ�pI�5�s+�F����{�i>J=�}o��;K�TI��T5�5bzwg��H葆q�q����7�)ɮ�ك�C�+?V�2�r��(��ߗ��3Ȅܚĥ��� _DV�?E3	q�[�}ǴZ��,'{Ug�v�N��)��'�S\���U�H|�Ǔ:�?����9{7G���+֓��Y#iƨ�q] YC<��o��Z�/(�A�7�!�7�/�X�_7�%;*B��հ�A�p�p��5 &h��g�r��`߿��y��ޡ:�����K����*q ��a�M՚�p5�$�9�_DZ����o�S�ٍ��ɵC�y�)�$س�I�;�+���{5��\�ؕK4s���l�i�Q�D��M����-�>*u�T�<u묙�^g�a�������p'�3*��K\D�oC��Y<j��:�&��h���Z���w��cTI�3&����b' �V9IBE��4�8b��)p+�d(���U�S�Û���k�:�1�n1{o<��En�\�=M$���W�D�##G#�����YO�
ֽXڧQ�y�&\��LL�癆��d�����vK�Zw2�4)�3���HJ�
�C����= �✢����;dG'���Ju6f}:Ä�4x\\.��J�q���1����F�����V��ET
A�c�g�%*(qE����$-�Dd�ޮx�/{��I�*v­�u�^;�䏍f:�|��+�LY��������|5&�K����UG+j���C���*���&UD�/�M0��N������z�$�'�����?�o	�5�lR� wR&m�fn�D�p����{�m���	�} �MX�8!1ͮN*�2�y7 h�׺ΐ�,
:i�i6�TL'Ṁ�M�;C��@U!H:�镂�RJ񒢖�4��ԧ�3���xq�8�!�G$���T�F�|q����ϰ��	zq�,O�1`�Oy�����֠KU�Ry�@�(Y���e)`H�⌃Wm=M���i�y�x�K��-��q"�����X;����Z���&J�Yb�Q��Ǣs�R���}Z�˯=.a����X����x'�=M�Xn�>9lM��hm��b��(��ڻ�3�4h�P#"9�G�������]S�W�f��k<�	�.ش��$��ɱ�a�\;$b���/V�!N]��x!J����m�z�3|L8��h%�[��@��O���y��8�?g��ǀW�����	�����Zރh��W%uel2@C��T,p�땴Բ�o,��O\`�Z@F���t۫i�ц�y])˘��.1L�>S�4is��s���)Ůڴ�_�!t���V؜�<���=����~�IE՟��bb�Y��n�'��P�m�q�L5"f��(|���*-s��h{L��m��l��'yq8V�&oZ�u`�N��~��T����d=�f-Y�?�Cv+x�cٺ��v�PMv��Z����4��%.�d���3��4�z�y,�6j2���Z]Lݎ�>���{��$<�ֱ53zʶiF�*$/.��B�-�!��`�Eb���s��ar4~w����ب�Ӛ���&0��&��Qo8����/3f�>{���r��K�;�и�Y�pH���8C9Cv��ZYS�;�ȅ0z|y@��w"�&�a>��L���:^?���-@���1 yUѰ;ÕT��";� ����?ɢw<r)XJFy<�D$�m	?�r�[�$�<a����P�!o���,n�T�+�T����㞫�pHjQ7����5J��V��
4�����:	�i�N���f��ms"%&�U���"g��e���p�Q�H �3݈hBz�i�B�Z���%�|�/o��8�5t*��XN��zY��9�T�4�f�E3G�8� ���q��4����S)$r`RE%�?�����+��/�B��oL���B�l+J���p\O����`ex��3d��*�{���䌱��?ct`�]ܐ��o::\Mؒ{%Մ �!^�j��p|�| � ��-�
�c��;@�����/Pg�D��+�
"pr��1B����8�'[��d�.�쮒�#ō�B3bȧqW��|g����O��y` ��F��{�	�Ti�%=�<�67�}:��]Q��o��q�����A�B�;�=��Fj��z���?+q�1������@�'�����H ��˼pHH���^��;�fj� �x$,�°��i��+���<˫�����OΣ�j�PM`�Y�L@�!2~���r���0�y�2�Ǥ�$_k��
S���}L�R�O��{��C��%J)��d���[wU�֦_��6�h��į]lB���h���׬r\�CNQp4��p��u�`6Σ�<��Q�r5�B�1s�Y�~mTl���g�ӱ}]�t��R�c�<� �߉+�=[�԰ZP���;�d3�+��!��΄��4�8���-2�̈́�pUL|�o�w��r|���������t��N�o]A�~DQ�n��F�c����{A��N�A-0T���~��p�M�he��pd#�W�~4q=z8V��&��KTd>�M�u]�p�m���ד$q������̀I(בۘq4��;����tsB<���v���\���T��&���%����i@�8�<r&T�
U�}:��1(5"�'��`1�fA�B�v@�SH9�/��8�"c�d���A2g�Hv�3g�[���O�IG���ƥ�����������a���T�a�y+���ξIg"��&ۡ�do^�x(�F<v�Q�O���U�<S�1'T�%������E�7�/�������H�<p�H�������R��R1�V�`��U�8��V�q0�O�xS3��W�mN	����B�e��o��\��i�˥���h�Q��x}�����~;���\R�Z����۟�"�k��Jo�#E��uTH���)T&h�\���$EC��xr�2-[�	DzA2xu������r�e�5A��q�C����7]�H��'Jk8�b���C���u+T�	��(�:�W����,���2�h���?nu�Z� �Kb�*S3���"�F:N��(�@�E֔����J\ϳ����S�t.��Y��v\+I�l$��?N����d�����=�x�zs������pt��0?���jgJ4HÔ$�.���HN��\�am�� �W\�X���?��Υ�\��<?5�Tj�f˙>�[�B�e�zf���:�Xl˯�evT
�b ����I�Qi��c��4c/��"U_���V���<��)e�XU�`�1H=����vP ,;+O�Q�����Ʌ���)�b9�9���ħ"m?1�GA�^Ј�9�bM�RU'L��w�
�nH>��*�/ߔ(�h_;>���Pj���[���s2��D[�����,��f!	C_#V��SEeyl�3��#����5vA��q�#^�itY�-������������u�S��{F �`.���&_�]'�w�/� 3��,���.]���U�g�(A�$�B$"]�
��u����r[�J ���8G���d�)�ׯ��Ply\ķD]�UP�(���>x�Ø�v�G�_�/LS�M>S�K0NV��b��t�"zP��bu��G����s�I�T�v��dU�ϧn�	td���>�tXĻ��P#��qu�.��9c6߿Z��������������J2 �r�.g�4�z���L�q����bpC��|z����6���t��ናw����UzO���=Ih<)��;��?]�G���il<��)%uM^���s���f��h��q���R����n�Ҍ@(��u�]�;��TĲ���+� ���h�d l�����+ФR0V� ʅN�E��M�0a��3w7(�����pv�&�d*\�˹E~�Z�g��� ~{�dU=n{�c��5�*���-O��(s�e�J�v�MJ(�TO'�8����Kp����~�ҳK��on�ܥ}�z�W�	r,��9/���^�F���V�R�ƄnWUd�p���6���j��e�����Yg����bB[�8k��2��W��3;eۺ]}�q�]�E���V;���*ڪC�xA�fy�U�Y�S���kf��";��q��D����3m��׆�7��?��-c��}���ǘ����ꣂ{9䇇2clUC=	�|J�I:=�C��<��P+�4-�d�靠�l�V%�gd�u��
'/j�NEX�}�tt�m#�)�e^����R4�d�?G���]�� :9y���q��C�M�jșco�FS�Q��F!f��&py��t�Ek�>�}��Y��n��>V��Hȫ	O'�".���X){����id��S)�d8>��'�hwI0YB�u�������E#���^xϒ��#�)$w�Ke��=#�c��PK�ճ��@�"�g7���$���H(ŉJʌ�y HRn^vs�i�2]+�HF�YS&�/��F�C���t(qt�7���&!��M.�Z���B��V`;kb?���@D�~��Ń�c�b}��|[�\�\ȝ�ᡗR)1�M�)�%lH_s��1@��QV�4҇��|��n��A�����B�a��'(A�����h�4�B�ws(�����a+f%֓�(���".�.!Di�x�Y��2vL��=!���T�OG0�|_�a����Q�����#�*�e��{����B3,������~�v�QY��f"�g�*��?JAx/���j��vc�)��+I��#�߅WSR�f.ƛ3�|O٨ݬ��;���d�4�90r��b�p�a��'i��ؿJv5��ߧ�l>N�X�,���TW�[�~N|V�1��t���2������<~��]ojwtZE �����l���v�٢�Pj60�3�2 �L��d�nwE�-0�lo<~�U@`	ȉ���+���5�V�F��Ii�.M[+���BRp�
�F��疏̑?���r	m���3�'�r��)_��G�4�v�H!�J�!�k����r��I���̗P�Z��կ��'<p'��`n	�9&��9sg�J���0^Ɣ���_,\��q-����cǕ��L�A�扁�)y,۴�O�<�
���Jy!��������X!�^�B�&�/�Z7`����I.zA��g��vabϨ�8Jj!�A`���Y@b�KX2���r�}�ss�*��<�z�0ޑ�P^��۔�ӎ ���(Q.<�6t.nNƸ�R����5�$� ��7ox�i"�����K"�%t���:�]Թ����������sS�i	�
��[�8x�������s_W�Ӛvv��#�90�f ~�:bj�X��eWu�A<�����]~�"���rL��wU��q�J�߬r���-^#~-�t�͝O=)�蟋��K��t p�A�=�^��E�B�)�wW�g�m�a��w曋�ySX�U2r|���&��	��c?����(?Q�aZ��E�(�[��՞�2��Ȭi��t�?kG
�pZ��]�������.9���E�<�1`�&�`����G��w���b'lI
k���3T� pN!��� ��`�,��&\�&�TM�H	L8�-q }(��J)��~<zJC�UY[k�m��BD�ȽS��ؤ!�Uv{7n�?�%#)� �|W�[�cl7�[���7+/��:���O8�8����ƘQ��ca��������i���5? ^���[�$����4��;YX��KI �TQ�/c�U��6�=�L)DT��?I�2<<݌ �e��.��h��xF-���8���f����z�*x�6[�̃�g䜔�*#�Z!;�ѝ�)�m*�� �$]��ͥ0�B$�8����\T��D%��C�軾{)�S�O4uB�сkk^ՔQ�7.�?�n��y{-������k��w?K_/�q"��YV�|�Y'[�լn:۝�e�v}O[�z�B�������b��Y��m.��<�~�nF�X��P��\D���O��Nߊ�4���fs�ȍjrd�Ī�{IOf�/���]��gΏ��'�؊�*�}�lc1��'^�v�� m��@��z�E��}��c-V� �Ψ��d-�
'`u�b-
�nĉ�d(P|����� ~`���~��~���HVDì��B�+g{��x͞ǉ ����4�/�Y!�����*���HK5�g����{�W� G�r]�6c��}F����Wg9�����.۲�{\��� �� ��d�7�+��U�Z?�\.؎�Ӭ��n���g�M�υ6k�^տ�G܈��W���w(M8A��i>m莛uV��N���q�&�v[��\��7mtm�I�Z��F��tDc �^��5d�ѷQ�V�Hs���󰧵�w�9���(���x�oMڱ��״7�Q��pEN�������d(&��s�;y�S��T
jF�W#�U���P��"����~�;.����Ya7XL��P$����7��=�fw�t����q�X���ꭌ[��:f��K&�*G\y������9��ϲ��w2�xb��nґ���C�u��N�js6h@`��K���5�U0oz֦e݋��.����`Qs�B�ˉC� VJ���~���j�/;D03Nt�!�a-����2G�Ž����I}'1��T��{a�3/>ߑ�,9PGF�~�V~E:��}Fw��Ik�'|���K�*Ho98:�G���.%�̩�E�W6���A�%q�A`u�^�ɒMёm�-H�Y��� �y~�>�-�^x��k>{1��V]=�sv���ev����L����j�"��*�!��t�^07)�aξ�{:_ })�`�~�k��.%�Pa�����ؐ*���cgcWP�Uϧ�\7>�����JM$/J|s|�V�Zx�ygs�V�
\�w�	ߴ�g��4;/K�
r�Y�3V��do��������u�j ��3�T�O
���4.���QS��1W�⪷����� �y��#������L��@K������!i��B$vX�����RJï��iA���Y�����Gg@:�O,d��~P��q3��Ww�B�
��X�t�sX�A�?��ޯ�i�8|���7ya50!��n|p���)�W9vh�	ZQ��R���ҕ>t�:�\C��ա��y�+�It�!H�Jd�c�e��]�ݞ�<��rI�sؓC�N��m��dψ��$S�XM�BCF������/�5Ă�ߥw'��8�4�]f�D����\����e�=.1xDױ�f�"����r>�{��|����m"��v'�x�c)�,b$&�8��vW�8id83�B���?,as�bJ�����ovO]	M��a-/64�N{߰dȇ����of?m���+Cw@-��(�Ä�Ǖ����JJNBA)�d-�5�L8=��"��:�ܺ,��<���鼈m�/��gs�E��A��/�(6Cj��!3�����
;e��EĠ31ޮ������=Fp"��+g��n�TQ�׻�R��%?]�Y��M��o�8B��D�Q,%6O@�����>�[�;�'��ɪ/·:㓌�[Y<���C��ԵAe�$#���;�"Ejn��jL����T-���T�} ��Z�\����gC�2l@4������~�잓ڋ�V��9����u�����,{օ�bAB�Z�~����ݻm:|����ҿ���&��K��E�Ǔ�\�ŷ il����N��\���G�ϹQ���Gq&��m�R�9\��,դ]��k>N=�,�1��K����}䶻*2�Y��$�}8	�	���4��T�#�ݭ�G"�L�ehB�Cż+�K�~���8���}�͑ƾ���2G�U�۬��C���-RI
�F����������Ҳmㅗ�Zh1��V�2�F�'S�<K��������in�J͚BA١��jTe��)M<a(6JfǍ=p gk)���O��8�w3J�n�/�n��I먽���]�X^x�!\�y~�1��B��e2��-C�.@�����l��I����G1���:6�-,�n2��=h��9�(����I�׌�[�S����{��7FY���4ҥ��L"�6O_|�ݲ�.e�iH�:!8��>��RozZt����ܗ��V<�J�Z���x�(A�ɍ1�uˈ��|�Ӎo_9���D���^���D�T��T<n�j����h#m!��P~��^�<Z���-���$n:��H���� ��\��ך� ��[q�vQ����X��8�w[%�����ò�`@!
�f�ǀ��.��(N�!�-�un7B�#���|`�kh��`���V�3�� �����,�c�H:?!>/�ʇ����֯L���_F�}g�ǅ	T���ɌM?�3�`��� \Tj�B����
S��OJy0yM���?�cCu��3�1��Jۍ7�C�4v[.\ʡ�%�9�j���x
Ҋ�����wǻ�wr�p�>/y	��b�څ���+��˽n�_�t3miU�-�2�(���I:�Lisu�����-*Eڐ����@�9��;N�)��s�)�s�ɞ\�9�!(��	شkt0o��6M>
H�c��Q�e���k,�ӛ��H��K�{���?��~�]^�.W��#���Ջ�����I�5>o��d�����xPDZ��t\��d�gs&�zb�T`�>:V�aG��Ko��[��k����W� zi��I�+Q�k��>�Nn(���:�8�<0��f�M*�*���_�VE&���q�!"����=1a�����o�$�����+��w}������*֟����UY�[��}M6��-� ���]�^��&������X��l:
�w�m]P48)�nI.@����������s20�����c�l�:��*�V�I)3cs�z��=��@T@����m�p�YY��*DF��#&.��C�l��u�7(��چ���C���w��s�|5aٿ0/,cceai�p���/[ ��Q*��u��6ա���E\!��C�n&��������&�a��nwEŰUk��&"��zO���Vp�KZZ��4s����zHdt���d��s"dx�@�=<�D��Q|C�J|xTUI�G:�ʲ��bX�̕*�&�V8��
Zj���IG|u+;��x�Yh8�J���@ʎ8���}�!_��]��&D��ۻ|ܦ�c_��':�V� ���8��"U���ˁnV��k U8[_��B0�P��TJ��\_��6����}6X�����A�ɘ	ɺ�M+�A��i�������QH�A�h�1��/=�M��fo8��DFQ@�Cw-�%H4�Zz��Z�����)��|����+��x�Sr��~:�Cy�Q�}M��-���p���*cQLg�L���>Z�z�Z@V����@������U&��Ak������3X{�ɝ[�K�(,�Sb�X��D�)�}vZ�4EN�m%���	��p��0`�_�X =Һ�Ul�t�NbYa*c��fRy���G��rE�?Y>�&��$��R)<�mO�Cysޑ��$%4�1��,�x��"���b%�~���M\RF�a���x��%��"�Js0��˴4�9TQ�o�1�ִg�f�]�![�E
��v8�$��[�ל��7��Sr�A��7'�IUt����*��qS�p�?ߙ��T�^��h<B,������ꯀ�����5�Y)�����@�{��`|O�
:�}�ӫf�-��z��`���P8.��߿����]sp���$i���{ɿY ��GՖ�<�*�|����0�BeI7})���,����+@B��ݲ��C��@2��I�)ٝmLeHrWg?�%��cO�цMOW�k����a��ڲ?�]��5�P��s�品C��k��S���S�������$ϼQ�R�T!|q B<:�W{s�
R�S��&S�b��v��t�(Q,���-��׸��	��"�����A�q��i�;�;!B�A��9�^�W��)�ej���e\�]�x-����Q�y��ߏ�8ͻb	�7x�×:;�?��^"���a5����'�^K�!��ܶD-��a|KJ�������a������{���6r���Y�c
�*Ϊ�ߐ�+�Е#���'���.��|& �`K%�0��L� ��&dm���F�<�e��{��T�` ��U�y%���?����_�o�-$�q@�7ƍ�Θ��u��P�qgA�"��߽7f?7W��m`���N�ڜ��+r៱�֙tqqM��Ob��?}��\`�l�XH]��Ȼ���F(Ƅ�a ��4��
��'�츍[�u��P�z�|���?걁U�4��y���	E'��E�!�Jv'!T���,��*�Xr�r�"��e4\���ՉQ��(�D)y��t	��bL�^Q�搜4���7��k�a��T�8ܪ����G���>w���I�VW[׷�$��f�'���6����`I:?C��M���%k�+Ӊ�֒'D�\���&�h"��4=���ÕD����&F?��SnVb�@�#%mK�	��q���ul��7��Q���f��gc��#lݶ�^�I�r�TQ�E�!�_�VD���2�K�~l&ܾ��}�U!���	����-��R ��_���Qv�U�K�S 4��\s;���a�G�Eqb"#z�����A0L�<t&�$����J2ᴒ�qpw��d��TՆ��Ҽ�*�+�W����H(����+{��T����o�!�f�P�	��"2d痸�%=�e����O�����3de� � �\ҕ�%�S�Ah�$H��-�;����TĔk�a�� �0�F ٱO�d6��'�N��\�=U�
�_*jۮcʕ#��?����5���+��I�Kb�^Q�1�J�`����r����_�����u�7S%�r#v��F�:$ax���]�΢U�Y���Kx��>-�T��a�'��ɢt�#���/�i&�O6� C���_tAp�O������}�}~���z�����|��c-�`Ծrwyw�9��s�F�#~�=�Gl���_9���zCGQAt?]lKH��u�	uE�GI�s��j1ތ���p�BJ��G*a����i&Z���aꢧ-��yg�A]�qL �MYU����y�.2w���UH�G��Έn�����s��4��WB��c(3��S���<G�8y1��0s����f9�$@�$��I��}�
&��	�x�ں?w�@�tmiV�=C�P�Tph�Q��P2�b("���p'	���:!|Y��Q����=��d�YF�t��^�VXK�� ��"Ju���sv�ڋ�C������8���i�h�w:E����w$�{6rZn	���Ҙ+�7�"3t5�z?8�ftW o�}��q���
�;�>:�nCZ��m�$�d6�e�z���Ni&�2�Ż�bs9��h���y�v�i�ҝ39��"��^��j|W���+�& $�e�	L�@�=-��1eR��yEJ ��i�����\M�����*�Q�a����j�S�C/TP�l3P3Gz��||o�tP��Oe'���z�ߥ���Mc!����[�~դl;�XsɄQ��K?��o���g,�����H�E�"l��Q��8��Ok����}�94�jѮH
�̨}�t^g~�R��ȪS�z��-����as��?��	Ke��R��DÔ>"_��qz���d�7N´I���ս��P�I�L�8ar�{ܷ��d�K��W탙�i+j��|o�_�9��j/c��a�y�!>kj9-����FXy�H�0F�W"��v�f�Dx=�$������g�pB=�R��d�Zg��
�[�z�>%=������&��mR�b���)"��4Ln��yM�5�?i!�L]�*6wJ9.C�] k8I�I�H��W�Fs��<%Q�� ���͢iR����߿���$��'~�]2�kRG?w�K	�VnP�����/�):��>���4+�"g����R���S]"[�O]� �u:��!ڂQ��ꋎ9M�~��ᨬh�Z�y#^�d.����H������ٕm���<ao��]�z���}��V���k����}�D*�4��h���TD���O��h����&9|
_(i�O7��(lʠ�a�K�^rMj���W����	C���3'�ͬ����S�?�D\v��t���H����+D%�$
Y%s|r)e��Ax�ZPT�a~i���=������̻*�����@�4q-RJ~S �6D�&�� ���/k�}�C
h�nN�a;��X\��V���H��Tɇ.�s$z�����ꧺ]�{jW�Jⶬ;:ƶYc�m	YI)�C$��~��-1>���C��a�~�5	nZ%8Y=�ASָ9���W{�Nr�����������1E0�RJ���m,XE�� 
!�H�W.o�GQ%�Ggwe�{��GҾ��������XG��O��d��G�B�:H�i�۽ِ`l~L���L�
_p����R0]&�	(�g�9"P8׊�&��T�#fx(��ɐ<'����rq�����q)���S�-��6{�Pw�eK�<u�fE�o��Eh�Y�w)�t�G]r㋢���~��O���I��ra���/�O�A%-�|vп�o��3*9Ѐ~��Q��T#��_��g8�d�{Y��.��T�"Wt.�#J=�����9�9�D_�3G��_@b��D3(����X�j�-vdM���}���|G3w�备�֏h�@��_vn"e�y*xt�&���w��su��P��U��.�� 7<�fv�������5-���},[~g�By0�ыt�_�WB�g��(������Wi�o��3�Q�`/%u��s,�Ea�O��F�+�vz��wתfXY*�ZT�V[�4�>'f��ݧ9�F;����\�h��z���S����Q���L:O����v�<��@|Ϣ��c�(-�/L��}\���4� �-3��`�r<� �]�7S�
i�����)��I���5�/b�S��݁���
�n���I��%�����AgեG3�iy	*�X�p��Ts0+��J�E�C��)!#�O8帵��ȓ�t��㋶�R����,�p�oQX��������T�M��6�����@�,	�6E���^��Te~de_�h��kV����!'�a;V���|C+T�F��yj�,�'�i*�n��-_��<�uA�m�j^�^�u��c�Lo�U�",�z����Ҵ�|��[���^)U�' ���8&�T~���]���Y̄o*�����Yfi��(��k���r{��n
�h�ѡși���s[�gY��ئ{�(�v4���YҨDiL�f}ݾt272o,�q9Z�1��S�7�+b����UH׶�J_/��Jm������8���4�b�6�x��ai�8��+�\ߑ.a埅j���tƖ&\JG�(e)H�� �^�E�;��ږ`������=�Ƚ����n�KO�?@�H���a�)�<徤ʿZy��CFR����j>٢WX*�ZM��R*L[�=\�nIq�ίe{1N��z,NX�����qD8�)���q���Qɻ0�����wOk�RA`���q*�lb�l�kZ{ʫ4��t���h��|�f�PS��$���=��*���YۭC����b�0�y;HS{M ��Z�sVF3�[{gq��i1A�t��gE\�Y@5J�G�ih ��$2��+��C��4-9bq��3|�K��Tȿ�Z=ZJ`ՙ��@d�[m3���pq�m�4�r�PQ��B���4ߑ��#�]������5�'Vx�J�7�0���Lޙ��\���19i����+[������"�Ѩ�d�`7P,O�� ������7|�ډ4��V��Y�M��@�l���D�6��b)��s�$���N���~.9�}���~��ćnJ�6����,�`��1����J�3��
�۹�E�-^�w5u]�k��I*����ֹ�YΗ�T`�`�y�8 a¥�=���Y�����?|/���0��ŻS_�e������\�o��w�@Mi2/D���qY��4��j��� ��q6utF������u��mOO��t��L� G��nk��yt���E�C\в��s5%������Pg	m��
`o�7���[��g���?j�'��)+wi-�38۔�%}f�����f��������^ :G�p[ǝ�K4@G4��>b���&���y�Fb�a�n�;�d�%�˨�u�g�������e��~E�v��5�_�I��ޅ��+1���0��J��m�[�rNH0�ݚ�@Œ?d�>PS�����di�p\�@�(���9�N�����'���v^v��,|kI��-r�w
�rO]F�7c���>��޾��9��l�:�sI�}r���ws
���s�j+�΄�|:�tW�ϵT�����^I��gZ���Ne���]��f"(�aDǇ�?O��>P�tk��^(n��b���U�+�ڡ�?�Vڙ�Wf��K����z{��ʝ���d*�|�w?Zǵ��@'Oh�O��k:	[��ތX��`库����	�5N{����S���*�����Q��Dt�茏����y9kL�F �$��i����A�a��HDZ��z����']&�躧D��2q���U���������o��{R��}Ot'δ�o4�5��e�?��*,��Im�
�a>��'�3W-]5<O5LM��j�7�G$�*S׌gT�R�P��o�Sp�&QW;M�6�9{t���.�>g0I]�}�
F��O�4w�S�NH��?X�8"rG%�M���Z}i������cl���tt�>ꌍ���J�$�}����(�B��G,�,��T���n|d ��XT� ������2���x�z��5u-�>�B���X�ԧ3U&�}���r����$����?����v1A]�=ڇ��_9�7���[F5��q��h.�Fqja��}�R�+���M����2蔴��
jq�?VS*���8?L�������5����Ϫ�lț�]�~&4+9���2�(z>���Ϥ~h�Y�(���w�%K�~�rD1��QL!um���]�M�|�� գ٥�;YN����5�'��H]�� �A^˅c�%�2��w%gK)��v��XP�{<YҴں��}VzG���H���F��x���QG���{|������P���q�ion�LO:�/�c�s\����w��n��Q�̀���1��<��7IH9�2�X�@Y�cF'�C��~[�D�����*�B�#0ќ#v�nE�;k���D���]bn���q�V�+&���%ʤ����z58z����ԋBL��-�+/�Cp	"|�������]�-����+�g�7�T�i�10�p瞄ϛ�U�sٜvK�� �6I�)2%���N�Q_B� s��T��i(����L!� ���X6�|Z\���'HK�>�����O�����Y�.�K^֢UKy=�'u��zV��2��4|3�y�~8s���_A�#:��?ǛV���o�3�'��M�Х\k�R�~b�S.���$n�!�', 0d}	K�\�@�_�9�mO�`�})�)MuάyKJ A������+2BM�)�N8�#]�<�	~<'�Q�t�;	���"�{@ d���s�-��{�bF��g7/E*�1u�[��tmW�����vh��z=z�-#<)�:�6��א�3���,U�!R�By��b�ԯ&����D��Ԯ$@ ��\tܾ��Ba�i:G#Udщ�b��35�C��sŸF�sjHݡft�c8t���~E�3u6ëYϘ�b���u/�=�H���\zLс��!�WT�9�\o&��0f���Kр��kv���^�2�d`}u����9#�Og���/��
�9�ic~��������~�^�e�1~VH{�䨛"����A�m�d�Bkjs� Q�,W�E��D�4��|m|�����1����)�,�v�=�.8j��(��]Ǟ��lQI��.��� ؂�QU�v��[g����_F+��޳�¿p�~�=a��y���3���)`�ܮj��@�*\���� �ɾ��;�ϲ��*9WՔ(��qKg���Pl����%��X+kw;PD��.w���lW�dЙ���Q%�ΕSZ�� �sPJ�.�|����J�}��p8�VLUln�I���3S[[�����-h-�4!$ּ�����n��mkOB:	��'n������ͻ�:���|B����,݀sH��;�f7#NS���LI����i(�`�VeC���S)��g�w���e��Eg�>Z<#\݀]�s&O��Hd�����%��nB2����K�Ov��i�V������a��	�Y�f���0���?Ó/�K�$���/��>8CS���U̩Ǚ�̶s9#�e@H�ۀ�4q�\AKT [����?G����v�"}�O*-2h��_Y�P������r"�i ���l��vk�͓�A��eЊȊ�m�:�=��f��#M�YL��O2�GԷ�����R7�@���tk��km�V��w���7;A�������]!��OH2�Da(�Q�Ô�o-A�JM�}��!W��XL��mQ��$^T�R���gs���~ ���ܻgYr=�v��Ƃ(�upI��,c�<��i����}>��ĉ}>�?�>H^����fz٧- �ڄ*�%�����%� f�t�r������}muv�)b����QIB��<b��Q�{`��o1��#��l��X��W�4#L&�<�x������<�1f;l������vTeU�k��>)$�Ǆ����(�[:�����O�kJ�����1�s_yT�����`2G��/���K��x���F�7u�Lp��T[�>��ɵe=��|ˇ�w�O�m�g���v����!����b��c���}����(۰n������P��nɋdǥ�)cnI�a۳���ϙ��A6�[c#Fp?��� e�f��<QGl+��f;���\Hc�zT2I�	�[[���
?�q�A���qpxT�8�bj�n8GH���=c�EʍQJU�j?��T��k~��ӱ=dfH՚�mi	�f���nPn���S���$i|!�fLd��8n�߅Vu� 3���3�� ��m8���g��ɶT5.��j����U����ǭU(�`M7��#6�c�yL\:�d�j7�_����z�y)�66>�8�����8�K������^G�H��!�B�������S�j�s�ɿӪ0�!�(C�}dZ��Y���2�V��eC�Xa�����4P��t�؍Ч���T�����++�_B����	��H����IԄm��5 V.�Zj:�@BUz�3�D�)�c�+t�Ր#��ܩ�:+B�L4�pl&׮Xz�u3��a���Мn<J�pX�h�g�힣u�|�y�33D9�
rC/�������U[�ӣ�p�?��L�M��D��l'�#H�J���"/[0�t�4���b��,��b��+3;�K�)��3��qG,����_�L�!�PDv�S-ō�W����X^��3�0�_���d11���S�n���Hk���ݞ2@C����!�L���U%��:%��m�SA��23e��7��	�˴�U�W�o�rj��d�/B��M/p����g�#�r�1{�z���՘�X+�뜏=@��s�-W=�բd��m-��-W�u^Ѭ0���ſ�zi+�����i3�]���2w��XfP2��[��^bJi�Ь |�bw���8�Vs3�KHn���F/+�'�?QP��\X�w���b�dr�qq{���E{[�!_1��WЊ�*�\��"p����[��Ƚ۾�
�H�����B�3���'���Q7�[���ZP�Z�L���⧮ەw����wНy�pzNm0�0�_w�&Q�.U����	[Q ��`�tc�_�۬X��(а���Xw��n3u� M1�Y'"�QzVl%ݮ��iչ��T�W�b�\N�`I�2�CѦ|J��)���_�|�N�>�#ĩ�B>���(���c�ױ���)ݯ]a�&��rG=�WU+�h=�p�ϖ���*��_#�WSi��U��?������U]"�b������8�w0+�L�?_���ݗܽO!�D,2B}��A͆*��.fU�|��(��������w'���B����ޟ���z��h���`�4U�XfA���f`aH��J��􎅃�>'��WJ�'�c|9XI�:Ɖ��C�3P+�8[F��=��(A$8{#5Dh���V���74��q+��*ɓ�\9��|K���T3�xϓ�S�]UKh��_��b6���� 0O�Fp�uw�r�U���d����K��t8h3����B1����~�A����ڋ����֚L�����p���DVT��BŉN�Df�Y��uX���/MÌ-��i�Oi���bzIw��[xB��2#X��v�Y�N3��l2��ib*�_��&�2[~ې�[��ܻZlp,C&wQ�~M_oz�� Q�M�{;,=J��D;���<t������J�����G����y��q��LDճd�����`c��"�����R����"ʗ�:�Q����'U[hE��	+�J�e��R8��H�%\��p�?3��+�a2�Mô���(1sdq,�ES�!W�`��CU� ��"�� J;W;YW�)�Z𣋮��ډ����oǾe�mT���bk�yB Xg:�Q�=qjV�Y����Cp��Ƅ~���=R(L��ki�{���d� ��x'����e@���ǈ��-�}�������#C8G�?�\�u�*-���?����.��zY�-��	��ҋ�K-�?�>L���.�W�X��N:Z��!c��]�;�Os
�aR\T�ҝ|ݣ�˂a���+is��I2�P�u��a�u1��]�t+��d��	״P!��֫W3~��#/H�.���zG_}N�?���^�)���,�ȥ'w"����b����������q�}Y���WG�菭�i�5ij%�pziq]�b�u�NZ+�0c���Z��.o�TgtZd��� ^~*�U+������@�J�[y��T�ň\ ��~o~�?�����8ݟ���[�7����$���;XT�SWv�d��U)#N��!0�зo���ԃ���ŤTՀ� p�H�p{3���;��`�+��Q[�-_d��&	UTH�$ �_V�u�x[��	b�@j �����	[�z63n�Z��_R	���譾�B�a�g���oV���b��XI���sA�&E�r�O��qh\̷'YD�ő&!�I��tG��U!��@���Ob�!ӈ>����#D�G�������\��5D�a�:�h��^��or���6��q�B|d�-Ǻ�)�c��a��2L�
ˍ�H�m�L`A�a�;v��^�*�%�I��і>�-ώ�ߓ��u�ʣ�f�*��^��u�R�z����M�H����s�Aj���3Yf;=����9�[鳏5�3\(�Y�&>�C3�je�yIZlf_�?�{쭵��
Φ+��ɉ@?5v3�]x#�E�A�J̓]�����s:�jR��|k���akU��4�t߸��� ����jEz�����k������=�c��au5�w��ѳ�=~?x�g��c�	�a��$������kY�.y��b��i�L��,�ySZ��.�h�"̷�%a�1��"�b�vq��:Q�8�O	��f�ϴݟ�oax�.�8/ʀ���k'� rk:JI���a�mw�n[ܵ��5s�?tw����%Z:�W��/4�����P�9/��s�
$���yR��w����b2���r��c|�w�F�်!^cz����˶f����D��Gx��y�[s�N��06t<"Oߛ�����7 ����5M/�Eq�d�P���z��x��15a.!����d|�욧����=����[����\L('���W9��3D��_h@�G�F���ʶ����#T�yJvtkO�S��3�Rq��� �o���K
�.�!?1�Ĕ���"�{޽s�>���E>��,�]��	 �|_��+>�=�]��)Ii4�'��I4_Y��"�Ry��8"1�>��q�_k�a��t�8Ym,���*sڒ�U��|��U�#t��I7 2�2�&��Y�}�ýuv�+���mZثN�Fr�Z��{_�ϱ0�\{���.��]�X�/�Wd�E���H"Ԡ�9�ǾnĜ��q�t�wb ��DS?��dq�^F�b�j�V��˸����4�����!����%rI}yNR&�-�'-h��� G[��L0�߲g�����zYO$�}��lol�����:mr��!)˛_�)�����5�wc���:X�%��l��o�Jݬ52�F��j�e���x�1[YB7�7�Ĳ}���(W��y\�Dѭ-3�5o�S�ZΊȩx�Fzn�2~>�P�
�>3���=��aN{����R�DLb$��x����]��"�#�Ɇ�G��^��ǎ��=D�n�3sܣ����2w(���xL��tcE-���a�COs�B�#^���<S����a��Є�c�h�X*����X�'Z^cg`�2&�����}�=��^IQ�k�`����a��0HL9�b�S��֣8l�_��k �D@>!�u���l�f�Q������.��eD�!"�}[ԯ�߿ץ�Y��I�Ì�_�s��S~z�s-R�9���b�!��~�5�J&@1�M�d6+�YF�h(䇊d�$.�����p~^�A7'� +)��g9�Ab�=�>A>�ڝJ���WN8�r��d��~0���dxh�6�?\�r��1@iq�nq�����������t'��Zn�3�\���dr}�㖔g׵O4R�h�9����X�f���>��:/�=�J,\�<���f�q�3�҈�B|�_����rʠ�4}�9��?�|ua|vw�]��i~ FՋ����R�ɲ�q�o#u�[^;�|kQ�Ҟ�OW�4�ed�87�	\���� ���ځ>G˨Ĉn��i�D���Ax՘;w{"������ S�'��ƪ��4jd�-W2:�wq�/�7��8�t�0��g1Tf�R��w +��#����l�Rˏ�p�(10%��'�bY���/f�9K�f5P�6+�Ś=�F���ǰa�wt~|���3�)�0f3\�IϾ�,)�	����>$C�nP��nR堨e�w!��b�>��``��J�mc$�H��B���%"a�i�	4�u� �S����D<����)�����<�����?I�&�sr^�tH
aE��.�cX'y\���:��7qٿ���h��;�p���<�Z�P��f��a����3f�Om�����7�aJ��K��^�TS�Q cl�'5�$�"��Yw��CtG��1��
)����
�;Vw�^m��"Z�����g/���5.����V����dQ����"(u���S�.U7��Q�80��[��耵,L�=��v�9��/k���<���#d-�;�)����w�k��%�������,L72��@�+">տ���oS1�#�@ۘ��;*���-FN�F�<��S:��)�dK�U,�@�"�m�-�%��2��l]%򟁊'����� S��M*AN�b�+�� )zH�	�����@G2�݁6ۯx�~�d��v�<��^��_`"���r)�"�/]�ݖ��0�*�a����;��e+��\�� ������P*>a
�u:3(0�>�h��Cp�{n=˱����:�����������lga�cd6�u��k���bQ���HЋ�uQA�71�l��)�Oa�{�����L	Ⱦ�G3#_E�UJ,1Ŝ8$ �n`���]���;�#\�~
���yz;*�B�d��JX��}�'|w�#�KQ>�38�����_u�?k�胬U��vm��W��?k��>U�}�o=~�{.�%�@���O��2&@��ɥ$�2 �Fxs��+v��Y �si��]<U�,-H��� ��tX���?8��18aQ����7w̳���/��4Jt�~�Kl7��&[L�(��]�߅��7�z�>��F�����I����η�;��-@��3-�hnٗPr�g� �*$[ݺ� ��A_n\)j9g��=����S�]�j�k�,J�2�
G!��!��Ɂ�����_1�
�vP!Lh��MW�Z��*���qy鯳�d���|:�9��Ko��;�-��I��HDQo�ę ��۽k�yg���J���)�@���ͫWlW,��a4�J�F�Q�pqu��K~S����F֭�^˛���}��є#	z��4ݳ&UM��>��}�	��KE��l�N-�?l�68faX�Y��a�"�n�l�v�������&Y�nk��N�y�T;+{~K�Ǣ��9����^��S��k�4���f7�����i�ֲ
�[����d�Q��������g�X�n�St�
-�����8��xx��|-�mi]��i��R֎�F?ƘD>F�"d
2�-�U��͓�#���K1~�5I���r�a�����̲;�A�?ݵ�Wy��D�>`�->D�'���Gx�?��+�a�Z[�_R����=Rџ����<��^߱xr0�V$�V28D�1�$�!g��;E�^�=_9Z�`ew[H<��xF��Ҭ����dՆj�:X+�դ2�獊��%xN	)�k�܅:+h6g�I<,�rQ}�$/�pts��3�I�Ea�0��4ި>��,�c)�r�L�F%RIg�����Ā&��9�0�?�j:����mʔ����+�HL��x-�2�n`s����hIl4�N77�b <f����Յ�/x,�9@�_���cX��^�J2�$�N�N��%�C"]����k�������� ����,��o({�T����E2�H==�r`�w&�
����-6��|
�J�ȉf��5j�^_� ř�{��t�^��ӀTDw�O	�g��b���88��j?�8��(��Z�����>W$�R�RY��	���p�Z�l�S$ڠ~�&4ק]�A�[3����\���\�^��w�w�Cw�
{�R�G;g�쓥��T��!�%"�b
�����k#�$�CA-+� �!A�O|d�(��f�~�f@jLu�s֥�(�ᶬ�k���Qf����]=W���K9���y�"��fJ�mL�݄������wʬ���ѵ����M}���2�;�嗂g\*>�+1�ull7��e�iAe��Ict
�������P+��0Ky|G��=xJ	�����G���h:���t.�
a��vZ����W�afq�0�6����Þ�8�
�r�v���" g�6��g�u&�q�P�p��qI��~�[�W���f����f�Z[��n� ����H������i��������B�e�M�-I��S�/8p|bb�!���CY*���Ņ�P.Hm�YX-�o�5}������y��1����z	�N�zGfU�����\���O��dA,<����X�~��vB�J���#�d0���.g{"KL�w��!���>D�!��>�&�JX;T�v]��#{M��4���_�ƍ���V|K V	_���2�y�Z�,�݆��Y_���	�JYL��g-V}g��z�?f�{��42�Nj'%�	RN~-Z��Іpm�J������O����El�1�6�s@�����hw&=0��ey�X~U�FOؑp~
��Ė��'�ӆ��1*��>ތE}{�8VW�B�t�o��5��P�lؙ�UHDh&���:wnڞ7Z���w\7��|L�nG�F��.��Q�"n]p^��Ē��G7��Ȏ���;+�4db?���;�B�7c������"�K)�UQh����l�"}�۶��:ҫ3�\g�r?%�9Gv�ޔ���C�^��'�K�ڝ���F�2�=���z���RvE&�?�g�>��Y�x/WK��t¸��k[�[��&�x�p�XH0}N�!�ZϹm���v�@��<�&|��~p�}�悑�K	��}���1>e�z�L�%8u)*�]H毣q���p�ö:Eg��bX���&"8�r���$����(�w�&X���mB8c�����~7��R���9�aޗ�\a�}� �9���Y(&�Ћ�O���( �����23p�h��A�.�
�#}r�Z	9�0�}PU�b��|��f
�9�uw�O�5[j#��q+D[s�NL��ԞL��h�n�V��W��r��%z-���ڷ���������Ӑ�& ������DU��@�M���.P[Xn�����ؖ��b1�pl�R<�׆�c���`��$��S}M��A�>��۩��k�ɥ[��/�WK�n�hrˍ������,f��g�0<��)�dp��!��;�+Bn @���1Ae��w�A��/��Q)S��`��*01>0YnV0 y��i��lS@'�:l��72�C��ܴ�K8�]8�∩�)aǀ���I[A�w5����b��X���%Z�#�կ�e�P�\2�t�\�{KG|.!��6���s�"�aA���sSW����Sړ.}��^D6�k�$^n_�f�5�-m���.�=Z�"�鈾��d�K�;i_bX}���UH�D�|B�7��y�*���$KY,����y���vG�k��4z�d��� ?N���դ�u�XR��k�{����K��C͜�:a?������k��/��ï�DG�v��)�I�5Q�!l��t,�����)�gK��<f;q'r~m��t����Kôͯ�)V�k(�h��� H�ύ��f��(%-�������[�᫼'�~O-��y�Uڊܥ9(̖��=.{^�:-���`�U�r/��Ѐ����`���_��r���rhp�R9q�]~�>�y$�����4�*�$*=g���`����K�:/��#oU�褙o8`�r@T����֥��'�~M'ZQ4P��}a�e� �G�%�l���	0oD#d�ѹ|���o=��q�E9߰�c�."�90�����J�i�	L{1\�'v�E�%C��xO"���xh4��s`t�
鉦�@=�3�����Oܼ�r�d��J��$L>��[6:������v!�4X�#�k%��"=>���Bֻ��Eב�O0=��9�a#���$�+���E[��ds�}�i�,]��#�D&'_������+][V	9cL�����O>"p�ɖ��#n�K�F�M
fY�N�~�@�z������d��oe���}��y51����7�R�9ai �^��<Np>N�3X��K�(�(�\����Q/f[d�N=��[��ڣ�NF5�rZ?M���|��!�\zE�����P�`Z ��m�t<�ryrif��Vz��Uk��� �Z����l4��� !���Ha����{�yz��ߙ�ˀ��G5��i����� ���"�izm��
��d���\�&	���c3&��?D���G��ylX
����s�^rÓ��#*�|�9���җ��hZ��t:>aL.��^J]��7�7�Ms���* �l�F��y� ?�X��
��=��?���Ea��o�vm:����OC<�� �E��]֝6����	[�6,Gr�O�	�_������ly�#�g֢FL�V}}VY6F8������A)QJ�FJ�����Ҹ�Y�#�=�@q�mтŀ���Z�H�6DUQ��,^7���?��Q#8�� ����P5?О���,�G�=Up�	7vo�ĩ��̌x&�P}���r|<8�,��G1V�!�9�4�� ��ƭ^�s�h��%U�]��룜����"��vʎ3�]� �CĨ^Z��3�R9h�
E�b�	��'��|V�:����";%*�g�GtbAA+����3����� 4�y�\�(qᮆ��[DYR�������,n''�f�u�q����Ly�8Ѱ#H��y�)���xV�~���Q�0fb4����4~�m{��tL��q��'��<���t5}@]b',�*Q�Kl��ֹ�2��"���u��D�`��U���):���M=j�73�9f��Ex�@��AXA(�ak�q8ݦ��+{3W���⾜��O��uBncsä���h�:�҂���]�?��>l���nګM�fB�{�,��6�i����K�c(Yy}>E���a%D��ٙ�P1�/��o7�����ާ�s╗5	;�r�����bbg�!�
6�-_��\�x��w���J9vsnv��V��s�X9����K���{k�=���6.�QkXD�"%��MI6���y�1�ᇸ��7!�������
DG:b�w��RҰl�R}��B�2��Ա��Xn��w����_�	�鼟�j��B$�qs�w�n��]��O�}�7}�Er�ʘ����B���x4�w��e�����'ZԥL9�0�	�c�<8��P�u	��'��%�ĺË�*`.�B+�cl{�Z�ܱ��;���ޏ�Vo�U�	�6[B��0n#1B���,�W`n�c?�L���o���)��{�p�Y��M]5�?�*v���#P.����n�n1����
HW�p�P�٪x�Hf��[䒮����_����Gs�����w�˭�'��Kʮ��>�\FOI�Wz=��m�B�^�Z��>��#��O� ,�rs`�'A�t�,�p�W�x������T߾.e1�7d�+O�~�C�� �[q�m�g8%�s	\��y��D���P��'wW� q����AZ�v�[��C[ti�~I�>[=Jau	�y���=��ٕuE���n�&a7�t6-?tO�./��a�я��'4��ͻ�D]3Iaͻ���Yhh��j�b�>_����ÓD�[����$qh�NV����&��'��!a4�6�F> y�Ţ�V\p��zg=�u�����>_��w�����n��˝y�y��{c��ǈʆ��Y$rs+��+~Թ�)|!#�y�Gk�O�%��@|I�(	%9��T zG�vROP��:���q?v_�n�%)�k�ݧ,����{���b�m��2��P��@u:�-�_��Nh�س,*��I�Z�۱{����͊��*T��(�̃("��H�Y2�����v(	�]=���JG��6j�����A�M4��?�A �)7�܇��8�����5�mp��8�����g9JJ����:�:̸f���paV��諤�w��^]����㥼y������T!3K��-� r7�I����S���$�[����a�0�:��@�"��]� �'�k4�C�Y=Զ�������V��~t�0��#�I��;�}�S�B~@���U�ӱ"��V<e��	���L�QM�ia %����$c�q_�q�<���֥�Ey�Y:��N�>Ǫ	�$��J/�p���&�p0��"z�z>ݿKfK�X򔖌���vb!)O��B��D�����$H5���xi��s��H��������K�N�W��^�SA���.Y�H#�y�����l�|�#o��@�s�>�s�*�*]ܚz�K)�&��Js�Z(_�;�KHR�؂�S���d�LE'[] DXg��E��:�\0���V~���&��I�UO}��nY��RUf��Ѡa��̂{_t�J�֝1@	��x�h��=�/N.��~N�5�+<����CT��ؐ7��U��N��W&�K�u��ꘛ9���ǝ�v���� \/X�U1=��;��I��>ߝy�Jq�'��`���UM+}�q�񢬦)~#�|S|QM�����K�[�g���M9ĳ}sV���l�ۨ�\�so#/�d��,9��ʩ�#P�1��=�I���T:l��9��eU���kL"�&���*EE���U���hpf��Rռ,�����z���G忚�L5M��bUv��w�Z���)u�pKL��4e�o^=7E8�&��`L�jn�{򰛻_W �Mx�ԛ՞�z�� /��Ͱҙd�ŭTE��l���͍a��Ԣ^����+i�ҫ8��܂��2Ul���;<��(3� �~�ʩ[��:w��0��|��]���&u骇����gk�'�����ndKݲǮq�ϔ�d��e�h�+K�\�W%�Vv�����|j���N������������d�/�V�i(�O`����'� ���z�c!.k�E��
�$�!ޝ��;��*�+�-����O:<�*;o.uU�-�P��<^�ي�^�h�$�~�����u{a
�A���w���&z�v��wCc�M����zCMf�Po5�C`{%r0������ǏɀØ�
�lH���2Q|Wվ�J���~*QW��f.`�q�M*0��#CiƱE���vPA6a�&&���i���~��o�����7Ao�*�����@uN���Zُ�<M�eYU�}�������8�Qh��Y>���C.0����'�QՋ�1X�C�rU�F��v%���xE&dP����w����ɋi?�
�@�e�j&��(b�6T `����yF���oI�*~-��[��Xlcp1��u��qT�8�n�=��� ���,�o�毲���������Ծ���5h񼁢��>2�_�(����`Lx�X�����Q{:{��HN`� j��^60�W���������b�@�"���		�6�'"�d<�2��� ^���[��� ���	d���疢�.-HY����$��+�4�;��h4
�I�Z�]����ǩ���6?�!��ؗ[^FP ���{�IA��h[�8�;O�F��V�m�jh��>��E�cV��7@C��vA�ݥ5'�vL+1�'���rEf���M�bb�ᙦP{Śj�)<ͥ�0��V��>vAX��X\��JRQ澐Rs�i�pY���VfB?���!�=*naw�R�e�8-/��T���:�K�-5��y�i暍�����]�1j���	��KsF�>��T���6́n�P#��	�ф�ଠ0l��W�,�b�L�R����������ZZ#�8ʭ~ѐ,\l~��`6�����:�;vANO�|��Xb�e�ࣲŉ��~ha���,ȫV�TP
�_���f,X��[�7l�K´���u�&�?�r����]��$�ۘɥ�~� "u��MR�"�	U�*�	�G	���U�=����̨��)�g���0f俇�H�{��ΐtX�Gc��#��H �Gq8J�t��e6PY�g�/�����*bS��InTᜂ�K������CK���T��_r�������`]v�d��n|EÃf�2њ+����;-�jH����ΫK~>�]P�S8������^��¨~/���k8�SD����d����-쐅J/1s��%a�Lbr��͜OTs 
ŇϓK��2��M΁<!1���6X�G_�] �.�+�����Ѱf��L���i��)�z�&�z���#�}����`3�x'Gt�YH�����5������25���,ߎ��d��v��L<��Y��2��t��sY�P�i��ƥ��s��.�0TH1Ȅ"s�FQ_N�K,��;�jA@��5{�%,�ÆO�=���p;؃�
)-<�&�IZ��m����u{_��&4L�Ԓ�+�T_\����	���-JRta׼�p���r}d��0V!���B��˰o�/������=%kԷFHt�^I�u�7C�d��!ʿ=�>Jt56}'\�y��%sW�S�M܊I!⦊x�:|���� �^�ʼ/��٭q(F��ki��1�"�xf8���%P��U�`*B��<&�����ݥ��.Ϝ)��iY~g��ڢy\K0OUp��d����G�G���;�����ę'5`���/;o,�I�8$(�?>�IV-�L^���kQ/8<T��;f�J��g����h$=].h�Ʊ�Z���j ێ?5E���O�Q���
T T�:���Gmrݏ*b�6�C���[r%8*G]�!y�3Q>�,����s���T��>8�����>!\X2����P[�Jk픕�o�oN�}j��4�Lx$��A���oDQK�D^'��VӒ
������[c��&r�X��ϋ~}P����xG��̱}�ɞ/0��q��n��r��n�w������l>E�A,���$��%w&�utr�U���m�ѐf,���im~ ~G)|m_9�����3Ʋ>�8�#�087l�P��4k����g7��>�Z�O��j4�,���⅌�����l2�YMw�3ePd��qY����XfHz�u��ms��]��C;��d�ЍE�j!]��~��(ȬT.~�Ţ��_���uH��KnM��y_�*}�$�c�e]j���v�vu�梅�
��ǭ<C2��毽f"�;�̕�H��
7-���j0oQ���Fx��H3O��ۮXʨ�-1��c�E=�Ybx?!5���^-����c��?�'�E��`c���������to��fWy8	⾸��&Un����d�d@�^P.�g��Yaձ��\w�2���p�g��hy�#�(����������׃� �h�?�rsj(]*�x^c�9�ܴ�S7����m����KXe�ϖ@3[�ӣ���\t�%ߡ�ԞMD�x��d-d��ܑ����v��Z1]���s�����'�N�7���`R;v�G�/O�����±�R����.н�i�c���}�x�s�)6��b�]�HL� ��1k[�����w�I�yE���\Y�����e����4��3^���]�}�|�͵�P�n�]��ҳ�^X�2��[Ռ����v.����
���\���N�kKۮ���#U�Ź��(O3N�jR#�6[ɡK&@��6�&��'��W�| B����(U�$7���)�д�fڭ~}yc�.����p��'�ǎR��p.ג�ym������s# G��4����O��B�sk������ �L�"t��� g��d����<Yf���F,-�{Oɧ�5wD#�ʹFZ�;���kB78�ّ�+�_`����b}�f�J���4]������|�2�u�;͋���}k��XH((�DN7gk�QR��F���=�~u3��zc�H��r�j>�j��/{i�+�@0m��N4�!4�Y��,T�+��S�>ȣ}����k�6���b$����ٴ���*�+���Ѣ��&�h��#��7=��R��p������hh8�����N�0�wʩe5 ���:$����|�J�A������m��Q�M�\j�[�+���"����#8�;Ƥ-h6���E<jI��Č�{D�_�|T:BV옄�4h]��C��ud��� ̘_�=��;��ir����=�P��0�)���O!�����3���0��En�k�H�t@�(R���3ypxp����W9�q�'-y�,C�bծ
��N��ka��K0��˧�IS�e���l��]U��z���#K������a!��/ոF:��~�ǜ[������,���Z�`"i�� �W�����sG���/��	A�N�\����ؠ%9����������XGQ1�g�ڎ'c�O~���(́��U�A=S��ʘ_X@a	L7��`z1Q�6�?+�/j�fE�͒�]��տ��]�ov�12;�s�#F��+ΫjW�3��3�;���9'�ɘ��� L��٨yg�!��-v����`ḎB'�ڛi�S��X7֬�1�CxVqY}�� ҈�_�� �3wM�M�E%�<N)�%����{E��̺w��/�0��z[NW�S�[<��K4�_�������0&gN��"��mU��|/ˀ:�jij��c�b�����KQK���t=#F�'�b��ۄ)`Z����VǱ��x1�����f�Z�>rT�P{^g���*����� �Pܰ��V��#]���c��$�O��^�Q$��ҍU���B ,�Q��QVSh�(Xb�wD��v8�V���ǰ���a���{�'����r����v����g���e !j�˖�T_DB���R�����i��>�I�E+�ɴ�6�����`�2n���2a~,��~ -)+� ��Z��z��^������چ�2g�܉W6%s�PF4�y�i�[w�#�Q��
��7��=�2j<��ș��,�@����������}�9� ��ioV����pS9��.�����]��rɀ`���Vt�yD�#��Tc)f�W	:�5���D�l᪼'��Nb��]�{����N�k�'Sa�r�6�ɶ�B"b����nb���t��:�TF��2~�%��W�;�S���+�~�j��;G�~�.�D��X2��XH}2B��uw7̉�,�N���u#$��l+�w��1�x"ԉ?��r��$��kv/KA��7�[�"��nI��Ap��r�-3�U�0�X���j�A3'ݲ�F��r�(KL����v�NU(I�¤I�YK*�\Y�B���{i:��6�N@x;���X�g�\��e��&�t��,;�tn�͵������ᚼ�����X{��d�q�3�jT�c�o�w���`�$����n��5Q�c���BC���9�ݛyR��Ŝ�c�ֲ��>�| ���_�0��KR��6xU��A^��.��o_W��G���B�CPF���Y*Zd)̋Tg�^����~�`��f�G��?�ɠra�Kp��}/��V%��Ir�E��	�I6x�M�WU��2�C?��L���[^�o��qK- ?��U��(��:���k�g�=��M�� :zx�nث���u�Ep�.О��n&��"&�L1��I��Z�mdbr��ʀs�<��r�u�8���3����)�qF��R�0y�����Ӈ�.�����Ϋm��b	��m����7�I$̺�Ś���vM�T�%��!Y�k�J�I1���M�]��X�d�O�92M����̻_��Z���W
$vU�N�&���N������D,M�d�N��������_lS�8��]M�>�3��3���M�����̀�i����),	��ޜ�x�@��έU'\��d�b���� �D�
�7�$��5��{�]��j�f0���aK�`&M��S�����^X?��*q	�R�R��J�4��(~!c9&�#_wD��֜|�R����n�uM�0_�c_>�ϥ=3&w��5����KI�����U��\W��x���s9�(q6��w*XK�m�ֆ��A���Ϗ�k����o(�̇=�mt�@�Ȭ��H��r�� d���cO:uM�t�g�(��b*�6�yD՝��:��b������t�xZ�d��|s`J��q���R���#���n�v+]�&�r�y����ʷ��t�כ޻M�����~י�n�5]�+�;'c��[��n�ЧF{ㄟ�����ArÁ�i,k�V�h�&Y�0P1��L�j$��54|W��ׂ�+������۶���\i�fEݨ�����)���L�N ރ~��Y]t��Ha�����6R��E��;==���6��U��.C���(���$K�P�����(�*~�;"n���PߠF`HN�NM瑏���d�~4;�����Bm���� ?�*���n_�f3���z��tyw�/?�h��b(�a�.&[���V�."7Xj��	���{���U|�� IQ��~p34{v��r�J��hC�3��kgv��U[ig��}NA�O#�-{����x��CS��e4����}�z�;"}� bf��C��5��
K�^��;-9Q��̋Jj��6
��ۖ�>~�K\l��b�0z~��OH���1\��`'�Wyl�p#����{#U�	x@M~����̰-6�a%P��!�NZR5x�����}�O�̴zlR�J4Yr["��m���>tUp7�m��,�:O`6y�.d0^qXN�왴&��Y_�v�������2t��Ӆsl�Of=y�4�yW`���!c�1p^'���^�y���0v�[�t���p�N����F��w�-%�`��)U�5��ҵv&?1j>h4����j�Ӵ9h���"�9�����X����EUQz�^�c�P7��Rū���c�j��b, ��>d� ���LUm�u�O�<Tg>����!I^Cȷ�i���KU�M�T8e(,+�`�h��@5��<à�q�:En�M2��Çc��r,[l 2�~W������{מ렯�����w|�g����qA7�|a,��I�E�-�(h[�:�+��t����*t��be;$Cgh��T�!ᮨ *g�GD���OK������jbN�δ��rPG������,e����X�W>�#w�VUѾ��<�Ԙ��>��z� ���6����y��Nf�0K2=�i^o_�|���E9�Y�v&�Bn�.e���q�n砖�I�p1�%	ΐ:���g�f~
4�N��%Yj��R�3�B��R�?�Z)A��(�"�j�t�;�F���:i��y�V�4�	*��y��s	�רqB׺hS�B�&K��L���e`�����_�x�B�cq��������]? q�yh��D ��?�o��L���D�=>�S>���#>�ӆ�:#�����_��%�#�4 ����<E�w�T$#sm#�z�I8�!{H2� S,�ڑ��  �4��y��4i��4�PN!J.�v�@*\N{����I������N���6٧�($|��q����0GX	9O���A�O�YA�~�GFj��{	�i�w����Nc��!u��ݕe˕Ɖ �Fѐ1ͮ�S�'6Kn�Ls7�+�)}z|�Ly�&\U�,A��?DԿͶfC�6�~_��N��9���x��EO��X����Z�16��=�4"��u�\9�I��03��bt\G����zi�L^v1%�:mv9��� �#�jTH9|��v�u�lIB��� w��(N�ݦ�̹�ĩ���x^�Y��ᨉ�!�{r��y:f�x7�Ce0zqP<	�mj��j�N7L�8T:BL��Ag���7�^�q %�/������ڻ��z�������zN����e�,��8T$7����U�z�ڱ*�WoR��?m!R�%��ž>X�$v�Tv�(�~>&M�ezV�C%�>���?��;T�|,t9��O�6�#'�F����D�/ɚ܏���ûu�
���p��2)J�{e��4�>Ly���Î��i���I&3<xcn��%��o�.�*3,�>�X�)��b;���2#Er6��:96�Lvÿ��lXĻ��+��V�+,����ҳX�s��|�<�ř\�};;�Kdlg�6ٶ��>�B�t�珈�e�A/�g�kc���^n�X����"�Y�^�Y��0���h�=YD�X~��c �|r��_$W�ϽCc��ej�&�x�E����/
��?j�>yǮ�nH�1�@�ʅ��#��7��_cK��:�M.�,���&{`��>�>6aKU��-�_��/>i�����!�S�8��_��;2��� ��Py�h�,X@��d�/'��@�QE �j�9���=��WT�-Ö8�,aZS����+f�v_�3qJ)�U6��D���4�#�������\��4�db�����n�g;V&�.�}Q�s;Ƨjo1e���'�܇	� Bl������5���C�@V�� �
����/�8�@qn"�~b�Ʈ�N����t�g��'���ٜڜ�%zi�2I�Eem�wG%��5��J��@1��������)��WCYf����ͱ���Rf/,���a��*Ra����<H����NȥS�hL{�AB��ܻ֚쾉����l�j:^a�]�PpAq����Ǧz˓~�6w�_{?U#��l0�(X��S�NJ�5�	}���e���̷eoQc�Z�W3΄��D̓����A���j�HD���P�Ԁ�9����0?>�cd�(�=� �n쀹�o�RJT>\��9��//@5,;���OG�E���v*]�*0yl���\�G�J�Z�@π6�[U��w?bSi:��e���~�5���<���I�n$�O�[�%u�4H��nQ-��b�8��;��Ļ����)R����Y@ߝۧ��D��1T,+�����	z���r��‰�X�u���rۿV�� ��O�|��>�;�*���3C��~�*���f�=����D���ò���[�Z�������RmE`�+�g=�
#��]^�.�H1z��S�Ku�O���LO*���	h�
-y��WUk���ݖ�gI��'p��S80ɧ6=;*�r���G�C^s�Q`�2>���)Σ:F'�� ������SS�������|R������"lU% ����ԭ���∦���v����s�Qk�4���jM��t?�S���/n��J2���	�?��`؛�u�?w9"�M���am͈hҪ��C1d�ާ�.�b6��D,Xe�C�i���y3�G���d��JY}���T<CGpT�J`�|�y/]����Cn+�a�(�2�VĪU��,�V��!�1�&���*���<axH���4�h���8C�z��8��} ۰xL�ΓwW1���x;οܗ@���W	0j�:Y���
�����gҐl�F���i�#�v�ظ3V1�d�����?$��N��:���mA�/���K�-Gd?.�5"jK�;�D������^��e��]�!7�Ϥ{��$��h(3�0�4���z�Ā���$KRb��O�M�쐍,j��|4CE�<�⢣. ��
��_�J0����s��%�{�Ќo��_�_�(L�4�����/�>7W*�?��g} [Q��DYV,�>c����ȸl�9�
!�C����SݓZ�t�0 �Vn\$&���w��BYM�(�?�Zo��:79����_��/cGg#	Y�*h}$��k_���'w�V�I�a���퐄��Xk.G4��Cԙ"�<�y�9El?�DߝLȌ��T�RE��v���$���~���k�
$Kk�~�2�˪��U������i4���_�;�6��-�`D� L�w`P��bN{�C�x�ڍ�,[τ!��_&H��H;e�Eg���%'-�Rv8��N�':�<��iL��īo�V*-i�'܎����!�[�c��}�B���-JLc�]I���1L7����<W/���ݵ��Qi n.���M�QG��a�_w-��ז���9������W�]��*  Œ�)0�,ώ,�c�d�lGאVʥ������h�b�������o+������D�ۨ�+�Ĉ�Ai{~��pV���������嚈��v+=�K�V6l���K�wT���b��x:kf���\X��Do�&�Zڪ?[c	,$w���N���Us�c	$xE*X���P�_2�H:��Q���C&Qt�0v��v%Y�4RJb�4i�^��꼫~|����A�qB4�F����΀���V��ߢfy-����M0K�f��C#��qQJaK
�	]'P�ob1Ԧ	.|�qhF�w��J��dnJ�x{�D;06<y�8v��r�(kؤ%�O2�A�)(r�=����.�hI�����̏"��ׯk�I�!t�zVf����Ł}~TɕO���' ��!��!#�y!���������K�+Y\�30u���5��
Oɐ�3���1��.��i�X7���^�i�+��^�g�<[�ZU\`}�	�Uby��8sG:��X{�qm��|�n���3ˊ4��{U���{l���=��.�O��+a[P�rC�Q"|�f4n�f�bv� E4��}!n�7��0z�J�r����,�>5b�V~����Mo�FĦ*K9׏-����e��:��Y-��1�D���2���2n�*}9b�U�^xЧv��Q�D�P�Ò����倨��V���-���M㶓Ԫ6���$u-l|p�0��d'�. ����/��K*�wF�A� ��~n0y���k�՟��w!a7�)��v-��e�.8���0�C¬ޗ�tF�M��h3���i��#��<Q����Μ)*`������4�K�%5D7�ɝeo%�YXZ��,I��MJT~�yW�r��z��xlj��R��_f�5��Ar����j���U�=�6k��Qq������!30w�� ˀ�g��M��'ŎL�\�����[�d��7Ն����t�10M�wv�l���<�W��J:�jCŽ�lbΙGU2���,�w���_�a���n�7�������P���VK��a��lbL��4�W4���E��oX?��tt"�*f�r�	�8J�*�x��6�XޓF`N��|�g$\��u�mO��gv'K �n���!�l�
"~�Z&��bTE�-���n�����A]�N]� ����Alz�U��7xfI]n�K.��A�r��N�嫑�8����d�s"K��a�A��Vz�Z2۰û�d�wjE�c �I&V�*1�i��3�7�s��g˶0դ>��uN��N� ;JR�.C����jt7p�������o$5\�q��∴�o��;*l�`Z������J9�����}7$���#���T�r��_
ύ�a~�ё�.�W�f^��{h�ңt���e����$C�K��^�.��`N��!zpL��~�oy����%3�H�X`&:dC�k�F��x�=���z_g� ��?�KU�Ұ�گ��Ê�v)M?r�rʂ�A��B�UF��A|���x�W���okP����T�Kr	2n�j��	�D_ʒ2�a��@�p��@Du'�H"O�{�u��B{�oQӢ�v ��h�	ox;Tٚ�1|�m�d��i<��	�^�Ѹ�@>_
�ݘ6}�}-fO�_-�i�D%��ө�J�f����<�_Ʀ{p�|������{t��[W�\��+��XG�	��G|*�8q��yw:ۇ;�'E�o;v7g��p$ (9Ҳv쭢�ק���l�{���z|��,�Yu6|�M} ��4$�����r-��}J>PI����+ڙ ��H��mI�.cT��*�6�B�Σ,^?r�+����� *���sM���?�<���ڐ����.ۊ���%��nH1~���	;��oQ�q��ϡ���5��n�G� ��4̃��1��3-���}^��}_Ξ��[���b#��gJ-k?\q����K9�n�^���>�F����Ff~��-�������h�&r�Y��)2���1�|�Ә;N�e�Z�����~��d)�;V��O�9Ojc'Q!��OIO;(f>)A�wlO��������0yv$�+u
�m48O�v�z�L���+i#�-?lz�$.��l��h����+zN �R�:/ٸɸ�q]�z��>����,���Bɛn��@��h��ߏ�xh��pT��4��f��&����d���aj�vC,$�3��4����gkܽ��ʱND�//�I�G)F��,oLC[lg����[�����߅�g�O�(�jK� q?�9�a˧�����e��U��T'ۦ/�#&�/ZB����~��MC���ANV�I��G�)K��Mѓ�6��9qx��ǒƄ��W��!}���ԖVn��%���-ߗ�8��iMn])��P	�L�a%�~Ӄ���T�9	6�5�p7�.�3l��c�и���s��F�2���>�J�ĹZi�7�]�	W��:� �AU�J��a�{*?>(f�SjqSqa*�F�A�4ac3�a�����SҖm��h��J�����4�ŝ�:��,ZݽD���Mt�|�����	!#'�N9�M�R>�XpM��Қ1`y�~	Ʒ�t"F2�B�.���L���a?�#�ѐe�lUq�$��|1|XS)��3P�f+�#[�ـǯ���fJō�O(��u���g���^+�
�|�E����7��T`V\>1z�.ST��7��b�~o<vv�wڠP&wMq�_��{�Qc��o����I�F�g�W�[�C��ŋ(>�t��b�~�حK�Q��q��dS�k���^�	pG[�Cn�4f��1�N5�c���[�%Ꟗ�\b��L��{�/sU��I���{?{��5rP���̆��	�iM����՞�.x�%������w��rkv�`��{�����%����q�ܭ'�鯔����%��b�S.0�3�N�&4oJ��}�#�h��,	��U�m�K�b�f9&?mB�􃌏p��B�_����jEL]L���d�"�_��>m8�ZZ%ݹ�����f�k()�X�?�����*�$s&Ă�s�V�cRt�9��%G�brdI ���J�/��Tfg!.�
��	CCQ%XU�UR�^3���!R�o�)Hn'0����s��W��F��M��.9+��+�6c�p��~n��^�D�C�=Pz���ܴZ�X�M�V;	4 �8�T�QݐZG�VHx��pgX� �k,<�^F"?������D�ʺR�Hr܊�pH��+b�4<�b�ժz��lB�W	��i���j�N��r��c^��׻����Yo����PM,N��(a����^Hrƫ7���;Q�dr�U�9lw�h��D
���p�G�i�q�L�t��~�)wf%~�m��<�_З��W":��f����Ig5EY�O���{n�����uqs���NX�!��=���L���$u�:�t39ho~��GI�Ϻ����XE;�K��^�)�()��0�B=Tc߁ƶ��Q��������3G\�7���!۾�gZT���S�S5�X4��Xj�5SB�z�*�m0>��fy�7���d�Suě��78_F=�$����9���V��9/.>��ق��ѱ�i,���r��q�&zӌ��L_�V�#�����~�M)cg	�#K��]��:�e��Gyt��EO"���S���T�̣�43l�� �;dEK�L����,8<�%�N��q��aJ���ܖ����N%/Cɀ��wA!O)Bs�db��؉e���޻2^�-hI�g���ֆ|��A=���R��E?7�ړG�ظ���̽V��+ )|�Ú����*����j����uK��
�>e����f�?e0��;t0pT�������-v�j���sl�k�5l]n��T0N����6>夠��W��zh���[_��W��rQ�(�G��3s��5�Xp��q9����a8buj^]��}�j����k6�ƣӗJ{�|J�Xk�E?	���N�MR�����L�ح�AA ��"؀�Iތ�@��DXKy�饪�:��cO��1î��/�2Y�J� �D����鱊�
x�9�ݭ�?5����I��Y�9�6��(P��w��u���E6�z�3��LD�;����~#��Н{¡z�Ae|�p���,��Y޻���6e�Aa�E�	�M��3ƣ��Q�7���%tF�r�'[,�0�U��2+�Fz���7�'6�b���NTӴ������!�5�28Lx����'� LJ䀘M@�Mc�� q����+9�F#���y�;x��3eE�ݺ��������D*?
���������\�1s��+���YO'��$)s/4TR���"Vh���Cז��vϩ^��C���޼������(r��T�����!`�I��3��x+��J;�au�yO�~%�$��RJgE�l��e�e-�p�����Q���|$��.���<.�|����<x[�3���@�a@��<������؂�ad��S͙&,���U�.� �J�5�=��lc�U�d�`¶ts�ʋ� �����Ч�?>��Z��6F�Z�U�{�,o�(�Y�j�ԁ��1�p�\���b�&�}��)� �u �2�#�! _�O����� ��h	�R�f��#J�J�D��a�s!��d���}F䏢*�5�7㣗rg�4���m]f)9ZL�	z9����$��X@kT���9�V~�)��[`R��#՟PP+l�S�7��9WV~�.��]�s���u�YM¸�5
I�؛�+)�h���I�-��Q�{��h���>W��`��e�n�w��Ǻ�����,�'{`�m�˄���N*�'�����x�6F�.����6���1�˭�o�H����wh�<��Ar��c�6�n�⒀��	�(��c�� �,{����T}��.�
�[pddڒi%C:�{,��i��mX�� �������E�wKo�(V	�.��bE��ltĕh�f�*������
��!�L����O=�� �ǎ�7��������'�{�U,X(?1`B�<]Kb�p#��^���ưР�8�q��iv)Ba����Dn7&#�8YtcJ	�F�AuӴ��B]n��>�� �	�F혉�P��W� �O�ݩo��@}��K�cOb��%�m*?�j'=j��krY��|� ���E�Uʺq*���t�N���B�D�aI4��F$my����^�zR��?f��KQܘ#�%���#� `O��!`-ه��Xt���;6	~�~�R����8���d���' S[N�	,��=2�/��
�([��xe���i����j��N\�/�,Vf��ߌ�[�X5Ai���?�N���Av��FA����`{��&C*T���N��`{����͊�k���gs��dm���Ӛ	^M��C�t��a�I)�=�3���/�:��w`�\D1E��*v�ͷ��Uv������׵���t
%�D��������sb4!H�B\�I�j���H�s�
�D�v��iɀ���������[̹�b�Z�U<S+��臨T�O������Đ�/+�*z;p�Mޜ)�w��բop��"]wRLj����	�ޱ|����RC�NW=1��z�C��df��>�WߑPuu�[t�oGQ��/$$%E�L_9��g�ʝŚlF1�4I��׵�)3/R�g���K�*�e�G�PxZlitkH-8��� �m�� \n�x+Ol�aD,vt��!;CŶ�e|�^Y�?�m�J����,:J��1��y0Z���.��z;\�WR6��Y���G\�L̾�6 ��	qn�+B[U�����r�6k{���И��K�����"��B���o''E�X��'����c3���;enty,�U�|�P{�_�Y�1	\) LEb>�&��~j߱[ipN�}���".����;��P���p��2������C~����}'ak��^B������S"N���m��1s8И��1��8�}Kdu�Q��=��k�vT5��(�Ґ��.�e�H���I�o@��f�=���{���{�<
�����YP���u�iPx�2V��������V�v���Ҡ��]\��(ᱎiP4˾�1��9��=�LJ+y�m�ޚ���:H��m�<B# �6q�O-j��bO�%2p���ѢrtM�����¤�"ڄ�={�/r'vY�J��}9��5�G@���6��r��g�y�C���pS7���铴��r���O�?�rƨ�(�3��A�����,�`��`Z�*�r�`�:4�sG�zL���1��?  �q��O>�әz�m�����矹qi��#�M�+�c�z�Ԡ:�3�� ��+,`Tw�Omx��@Lm�_��e�F=����^LAd^��RO4S�pxP�}��53��c�}�/�N�Ʀ��9O��Bu$���m!��]*�+��8�|KҞW�*���F�k,f+�6���c�sD(�y��2)�3G�g.К���\�
��eOmƥ\l؁'�-�z"˱?���dи�#�;,j��.�:�?��2�R,�tAb>C�9� Im`P�NVw��#�P�4]7�->~Ԕ9m�"��J,�_�)�������x �թjh�L2�=�����Ӿ|ܥM#�qVq��1��mM�哦Q�L2����Ш����Bl�pWҹ�7na�)���50��* ��d*���RJ0V'A�#՞s9�4�W��^ ������O��	s�I�&�� �������� ��N�Z	�����6�Zrigb��f���{Qf|D�	hS{��H�3v��=�� �G!%Z����Rei����N��`�7/��&�nCfM@+M)�7�`�*?��u�����6#��F>��R��u#�M@	-�3������B�Wϲ�H�'7C�I�{�Mds#��8:����"�M����t�λ}@?�OheW-��Q����#M(�pm�[��.���̢�^�Q�z^�s�=E�)h��P�;��b]ޜy���F�X��M�"�\,���6�)��Z�J���Tq̣W�	�S�#޾h-Q1�rG�E�w(���:����'2�+xU�lR6c)�זG��\�3��0h�����y��֧��6O�1�4 ������^�̡�>q{ 8Si�]N0���4���4��%.�,��u]�<�T�5V�,��ֺ߬�,<��K|�"�wJ��.�gP,Lk@�;FS�\e���6�i����UJ@��K�|�+
nZj.���x���w�/:1�صݓ7y�s���J�_��.�S� |fƳ�ߒ�{�C�����a��5[����d�#UUI�^LY��5ɡ,�p�d�f�L8X��bQ�& t�N}�|�(J�qM�:�/�?CgG!h����pn�D�q��]u>E7����nMQ����;�7u]��XL)�Un�[�����&�s�	�����ܠ�Eb���`M$N	N:�� �C��kM�r�fpT|T>��!]�ɵ7� �c�$��,��yvQ3���\4�z=̋v�:e�wk�N�b0@ܺ퓏�d��4E����F]#�� 	�!�y��H4]��2�3�_ u�3��au�}hW�*�^���2pJ����ɔ/D�I�F|:� #�Y}oI)-��s�q@�?V;;� jW�O���3�9�㑎��݂:4���2�V�P�0���'/���W��_CP�����`�Q���ɉ��7L��x��O��B�R�Ӵ�H��K���H��(G�5��.�Ky�K8(�LGEg�w	(Z7D��dꥴѕ�`�-!��sd�l�a�M�C����M�G���>S�Z��:ֺ��1u��J=��k:5���Ro���hԧS�?�]�(zT�ʛ�Xɓ���6�݂��w�Cf��d�tZ��b���v�EO��D�期	;Q�1.�)�ż;3`��c�0G∹���8�Ge%y�*���
�^{��5C���]>m;����	����:*qG\8�7O]"f�D�j�&�X~$A��Ϩ�P+����
��(|�ķ�xIQ��6�輓�Ȭe���V��>zs`�h'E�"�s�ؗ̈́xc����u^�B
�$��hQޱs�Ƅ^�)r�1<}�����N�m��U�@�5�稱�-O��p�{��VS{��lj0�Bo�(+h��
�Yq�U�2Fu���I��\�բ�l����6�G��V�K�m(����r
�����S���`��x���R�"�&�HN�b��d�B��H�l�'�2POb�諯�%/�W��}}�S�fA�M�W�ǎ�����b�3=�����w��zԖ���s
t�,�I�'�_��!?�l�Av|b衑f�$�=�{r�[Lu��k�<3��¨/���E�SqԨ㲖����k�K�zQ�>�#)�>�N���tL���6�9�O*��I�Ejaۢ����$9��J��tޒ��dB.�)+Ϩ!�����&����K�΅�Кf��uy�!6�YS(���f���&d_O�y�$����W3�G�ě6�#x���,��\�zWܘdI"�;��pM���;��k����h�&q'�l)j��#���	�S�<��G� �R��q��#+�#<:�+$˳�r�zJLt�4�2�g�>�(%�/Ֆ��d���y#�x�$��u���FԊB ��z1=gk��:x�1)�GR��J:<���M�uئ��.6xjg���2��v����(M��H�G�P�_���0�k��nҜ�8�Tz�>���3�{)�p��u^�g�������r����xD�7��E��]�}�K��{�F,Oq���{���~�U���Ԥ�]$N�[
\PsL#�#M�u��"�I�l��O߭�M�W%�c��z���-���#�D�{�-����B�L`��7�ø!k�?�ۆ/f�L�mR��ϥ��"�-&>R�~D������nX��_��JY�g��_od�1ƹ����	[Ot/�E���x"�V����e�%w��{Y����Ҝ���Ae�lE�p����@�řH��}t;,JA�������:#��k_��/*mi���^��I^j��t/�* �=�����i�`c	��}덄�1*��������I�uβ�;`�"�Z)��a�,fV���D)3��c����#�����3�^�HFf���6���-F����O�N�Z�:�mO�o�>G}�˝��V�%itd��r�:tId��0aՅ&��6/D��ǲ���UC5flJt�8�4*�WW4n�/Qp�]}�;�Cr���`�qS}��Ԉ7�M/�"��}$P@�}� a�%�]�6vԯ�Ԉ���t�˗�}�(����PgV� E��F/��mFioD.	�e���ǹ7�n<h�7��B�Z'�76�I���_�g��"b3l�a�~���ø��A$�u�Ey�n>�#����]c++$^���Ҁ4����"���c�ˍNo��*R���0k��pŴh
��]Ry��+^]�#�/�ы.A�\�)ځ�RSt���ʒA�N�[+~ϼ�F���&��z斥�Ђ�t!y*9�Vh�c����0�ԇ���n��#K���d�hr��@=�q��U�$Z�C3WAL�\dB0�6�ꛁ��2�gթ��F���d�d�B����6M��]f��(�)9�C	���O�/R��ęR�}z[�T�1rqY���H�j��k��N�i��	���P�茘���񮌋�>1� �Z5jo�F�AE�&��	@���y��[|�z�[����Y�X�2�mA�+q!���\�e�I\�����-�$q��x_��G ����Ǆ�W���~B�o�(q��F�)"��1G4����
1���^��]��9D��n�+����#:,�Ec
;�DӲ\]�N(1��OlIr�g�a��v3�+�W��+�������Ka���8Kt��-,
^�gTJR����'g�y��������dC@�v����)�a�[d���Z���T��cȼB�x:\���'��8�\����kγ���$(Y�䧒h�{�_IS"R�-��#����lU�n:�t�_���/�-Hj�n��2'�̌�����) TZ����o%{=Q���l�GK��7ں V�nZ��8mn�f�t��04�9W�,��2��1^Y�W!�'9K��)���g
X���$��;������\f�׆}�2�[?��T�v��=4�r�:��PBx�����t��|�N8� ˠ�� ���j���op9D̈́�?�c��V5���o�=VQ�U��,7-����PYˠ�z����V �D}\E�0�ĻS����L`�=���<2�����t~59ˍ�}��4/7rL�W'�2�}�E������x��sؽ�K�E4�����B2's䟐vFŢ{�>�G��'�!�؏���:Y]v��%(�a9"L��U���9�ow�R!��#����'�$��_�&+esZ x������v��Ac#�N�����Gr�	��`~͜tZ�M@a�Ĺ��㈿%%鄔"��F)$Ȩ7��[cLǮw���u9/� f��f����]Tiw���6o0p�-��'AD���.�-M8��q�W�rԖC�KVy㰎E��[ K拙�v�^I���~؛��x�|n�S�o)���"Jp�f�o��Z����iq�&�9P0j�D�m�_��Cy�J(�K�E��d��8��O��wM0���z}[$I$�_I��=}J*�����Qi1g�׀!t6r[��$~����+5U	Bq�X�j=358�Ϟu� 6�<���g���h���1�ľ	����<�ʍ��ki�/3p�������v&V��\�bb{?_�aS��{9���
�2ӷdd�����{i�.�h~ 'I�"�Xq��ި������FYG@D�#����k�)>���I�c����(%�UD}a��#�H�Oi�^Q]���̼tp�`��@R��pFNpNT��Aj��0�97Y�WW5��l9��t���X��(y$��~� ��Obl���&(ڣt�$��j�aV�,�hf�L.q6�����vG�2�l�L�����\뱲�GXF�$���:bܥ��:��Hʖ�<����
~�ĒSUï��;�FrB���p/>�"����
��9��2;���TA}U|�vʏB�ClQ���uYZ�Ü��-y֬޺��bHf� eB >e%q	Q�4��=���i?�<-{���Hö��?����<��ꌖa3<W�f5�i��t��Ć����k܍G��d��/2��^J�s�)���i@�buʚegRqo�}8x��{��@DR�Œ���+�X{=z�&1vy�������6y�ZD�i]��@�IE�8&AK4sX]�&��&�Ն��ݐ���b���]�+yl��F�m��p�$�C��闎5�qmg'�#�60Y��
FC��l��<���儝3�\+�?��ʜ�
_+�Ȣ*K_']`�� ���j���hr��z����B�:�Vg��Nc@(��"o/Ǡ��#�{�֌�����#��b�	~���PY.��ӡ���9���ʑ!yҎ�ש�����o�5`�wK�=|<�'�c��|�����HG��A�	k�N�lޤ�'l�S�o���ޥ�T@�@�#��$��Z���p(�
녤A�ш�9k>؆�+�ܿ����#WZ�y����e�|��<���'V�[z��|sɆ)�kr�5���Ś,	�
O��I��}���Y����)g��0A��dsH#M�,&s3���?��\����ED�a�p�쿶-,�:����Zf�`�(Sv�1�/s'b��ؐ��ۄ�즕k쥈�R7���y�&���{�oAO~���ݎ�GV|��3�!������LtsZ�Vlc�xH�8Xb`w��N�o%�Zu�Z���͝�*"��
b�CC�ϻ������`5Tz�oh���b�e��������1L݀�9]�����K]�0�k4���N#�C�JmxO�:����\#YN ��i��V~����an�J�+b�u&��H���r�O��U@@&~�g�V�g��.-YL3�v�)��&/DLzI]L��Z~�(A{����YD�XnF�2�[�����B����[
�G�Hl��w	,5^��g稑*OB�=?8g?VW�}TH���9dh'�;eC�Pk�����w��ϴkk��E�H2S��m����7���?��n�K���[0|��-�Һ��r��9� V�U�����x����4�DZ+r�ӷ0��o?5!�w�#�e��#ʱ|p�wd��4��[���y��i������h#�+�m� ���	�S<2B�sm�Y.6�w�K��|6j����is��$�Γ���#�?i�����RD=���2���2��M69��R�F"J��t�#o>��@�hx���z�4�#u�,�"��,���#k�1��X/���Kj�2���'��y����imKv���^ʵN;�h_N%�jBq���J�c,��r��/�y�3�>+[<�-�oz�m67����=
昗��m{���"%���}��+�렂I�����ˬ��=����'��b�αcD�e�	[�'�ڒy�<א	��+q��$U�F�lM\r�k,´'4��g����)o�/ijh�MZp�W���`n��s�b��p�O��M'�����Aձq�u�f쌛�����.��)�?�%��jeC�Ӫ�r ��]_��0+~���� �scI��0�=xV��6��?�7۠�7���?+R܉��@x�o���{q�;�Ir�jۍ��n�V��Se��ܯZ��={E�x".�{��W	3����=�H��~���"�
���1�*��G�����"}5Z7�L.d����2�@m?}�l}��"��:sK������wm�y�2�u���mv���j	5ZCi��.��~_�N깘��� 䰍ƒ�Ը��*�{^�t�קxb�{�Y�xs,�
�WĐ��sV��T��k��/F�.��ݶh���T�'�ZI���I����&t�����$͘	,)�.b�7<�o�ZO�`LB2�(ݟ�o�v}L�A5���~g��3��|�h��O*Y��fxi��Ǎ����0l�?�PO��d�b�H���f���\��=�r� �}Mc��<����xb�K�ꐏV�G���l���gz����%r#đ���qD&�_�/��c���Ӯ_��3�`�ySmF�s���)�V�����R���'N���ϗ��	Q�KsJ�M9D��w��.*���䴨9�L���fN���?�i6�K$m�1�@=�U�O�R~Gd�Ng&��n���'��e���c�4æ��a������%�B�E]����~�.��R�s�]�uֻbOe�Bh�:���w��c��$�Zޘ���e��իO�����㲜N��(�}�Z�� X��Y�S���M���B��J�۰۝|�+�$8�-���3����l�.-��Fou3��5�1X����n��6�'�~��|.m�F��gKH+���j�WU3OhV��K�dJ�ыL/т� u��ů dp-ܛ�v�<��.A�/�ǃ�j�"��Q#�����j"��'��������$�$3aÓ�$O�X�'^O���	�������nUS�9��to�;.Y��g�K�´�pN����Е�8�F_��m:��h��I��,��i��Q����=s�#&~������ � ���<�b��n�XyI>�q�W�	���"H�� _�� _��:إNB�jt�K�r�h��;�EP�zl7`s"��Ȋ-�x����yeݯ��ʻ�ö��p��s�IO<�Ĺ
/�
s���s��ځ+�Ӑ�"��v8yhi�?/6r���x���8���~Rp���l˾|XLR��q����BS�h��� �>Ƥ��V��Z��׵Fh�V������[��́h� � 6%��\�K��N���f�?��|.Eq���>�Ў*0�}��Q�󱁮�.�я����\������2q"i�w|y�PN_��t���ȼrʻj���x&�ȸ
��e�
i�a7�.6bS��t/X�뒔�s�hN�rdW��i(~H�Z�����"L�{n��R�:�p�pqb���_b�ts�q�I�a)s�_􎛨؅ۜ��a�u�j�6��NV�;���S�6!��XF�_u�W��"Ɏ�]�}ЊD]�	Z���}�H�u@Mv_ю�i ؁�|B2�c�&�`�L�(3<�@�Ag)�¦[�҇|X�������z�H� �L)� ��)g�������.L{D6����vʫwE�����/U�^P�]�F�?Qk?���ͧ6_T�S񽍺�$���1����Ш�F�3�@��Um*)�N�����!k�[��[�oV; �3�}n5	O��p�O�cY�ɟ�V8~WO6@�zo,>�=�{!K;)?�!��y|���hYB7�Gy{YGN6bi�C{1�fӰ�f[�c,B\◅6���$m&����_�<��"r5��vǯe��C����r*~�ʫ��RL=���{�O�=$�GW�gNR�њ��L__�?�N��aQ�D�l^!��O ˘6�?X-II�Jؿ�̊�:r�A�c�)y����4�y�>�́*��i~��%�}A����0��w� ��p9A�^����a�n�wr���\��	&)#釪#��yS���<��x���@��E�|���(Ut�)��Ϥ���Ɖ�8�`u\�612�p���k�& F��ad�v1R��k�����G�::����ˍ�*��}J�鯷����_c���x��|4յ�i��_	���{�@��tjE  &�J]Π�Zg	�W&]X�\@� n�nQ��*� 铷]h1�zVXDS�$�SRՆ('�)����)Ĩ��$7����_����Uʗ��\��0uX,�z/��Y�u�gOl�7p�P�͖M�S�����-uTD�S�?�ƣ�w�e�E��~!&9�9�b�h��]&w�*�$�w���n2�mT]������PL#v
���id,듂�S8��iݝ"VC��؏Ɏ�l�}X-m����,fc���>�⶟]ɠ�����M�� )�9��8Z�.��Zp7��h�{�k��_/�5�����gۄ�ן|5�c'������U^��M ��/s�����M�Sy
��=Oq'ו�b�l9�/� ��
Չ��q6��)p��S���_ZZ��������C6a�a$-��of�ߋ*I))7��]�zg���Gu���ѶYB����o�X�!NJ�{IaOf6dS��p�*K��~f�\K�|P 2�c��`�D��(�)��չ*�����-PƘj��p���Iubca�6?��#�e�����pŅ�����h��޵$�0���ae3y�IV�
�;�hU�!�Ī�]ץ��dj|c��7`��	p�F�%�C������J�@��d��V-���O��ɑ)J����+��y�X�UUW�A��b%�Vѵ�sm��!�h?�	��glJ��%h�p#�mv�A�f���#X	��M%�4�>��/#S���xX�A�`,�H� h�ا�v�rU���-|>e�@9�St։� ��e�QE�K�����|+�X|����k��GG�ה4Q'�y��8�.�n=;oR�ȁ����`� ��� ��&�j�<EX��g�&L�r&�F�
�Ɯ��0݅�g�v��\��n��gZ6h�}��l7ڛ���I�F�#��;?�/OE���tI �1�XrR�u͘�7�*�4W�����^�P� (6�N�E��V��X��A��:����q2c-�����4z�h�j���ݣ�8����C��Y2uw���'m�#
�7��2X�Ɩs����'Y�p�̴�w����f����Os�Qn�K��u�&,�D&�AD}K
��=����eOV�zK?/1j���*Õ&���|�4�������||����� o��+��@�`���߽�x2�{$�nr�/׍�nm��l*6!v{�{�*��BSAr�.�jVe�w����%������Or%io��s�U���s���0��i`�ؙ���Ԯ�۴^����O�sx��cy�h�]�m	b�䪏�׷]S�z8����3T~7WQmO.�b�j��ݔ2��x�C�'՚�3�ż\b��1Z:F�����'K�N
Z�+a���اK%� ����л(�G/U�U��-���q	��W�s�� �|�������A��+�
6Y�#'�ϲ��+�Y�0�;�-|8FܥF_ �K¶��GP��,��X�������AEb�qډ���E�P7���pP����8_��'�;o��2�s1�Q|��{� t�|L�;�	��Ro���\����)��_��hO�yZo��!�!�̒�f�I}Z�LGڡ}1t�N�~��?�a<@t����u�l��߼�5�������=5Y�*)o����Kn=f�+��VJ�>�1^,������/A�e��J�Ñ3$C�g��ؙR'!���y�Ԁ6�V}�[9u{0�t�FB6����7������}�BP��F�������{@<�@���<�����v�e	��Tx�jG�$��k0�)��k��jM�&.�d�G@Qa�|ݯ�z�1|��6{�6��`�t�_����|��^b\�4����CI�f� ����Ux����㷝fܲ��*Q_@XD����u>U�b?�J)Seg� u��E�������lTlH�w��'+[&?Ğ��F��D4��;lؿ��e�+�%��5a��:�2b�ۚo_'ߓ�L�����Go#�4�;���Y�,͚=4Ύ*���h$���s�]vm�ufHeib��|\�̞l��0����q1[�F��u�mU���l�J>��j�O���!���" ��$;�A���>����f����&���l=H�G���$Y"��W� �k#�;�61�R�zc爒��5b%ph�N"^Kɋ���k�诨J�ِ�R�R�v�&��8�.t��%,�}�9Y�wW@,����|N�\�Ou���~&���~��u�K�S���X��+b�sy=���%gU�� �����g��&��C`��N�p��OHL�8�lth���/����"*V����p���	w�Ճ0q�s� ��ւ�ޠ��πC�,ZW�i|��Z�j�"\�7p LmkiS��ݟn�O~��n>�A��2'\"VnoZs� ��	�B-��I��4�;2�)��H�� {h=f�;)ܞ]��/[��q �������8 wg���u�p�巶�?���]E�/����[��B�%��x^���/H7�F��)ş���x���+����YE�=����> �l�w�{�b��_�~o���F�޶v&��u9�#d�i.H��'S��ݽe$&<�څ�x%�Qg�ic�#?��T�&���
��A{}q�#Lb(�����b��9nP�-�G��� �7'Td��������]����bT�c���F��d	�!�c���;��:�.L�1[<��ڢCU�ST��9���q�ڮ�z>TME���$·_=B�P˰?���eW"��{No�ؘE[~M���N���	bL���Ͳ�ޔ$��K	�,c/��qzCN�A0�t�pd�z�-��p��/���-D�F���E#�Q�:�z.�P/�K^���,Dm�qYi��F�|��գq�ahj��_�-k�Q�ƛ7��p�E�H	Cl�Z�W`���'�m#_���o�������9�G|d�"�~f��;�@4��<6�z�[吟��[Ͼ��/�E1V"�'Za��w����U��@u.}-C.�~�����oV��F��F����ߏ.`��>�o�V@%���e�����K��&Ԫ/^g1;eY6��y�ͺ>
�q7�ވ�s�x���4�=R ��QxX��M��`�3��4:���ǉlX�s��������"���D��.��5g�=	'xz��Z���B\7��O2����k-h��p�Nrژ�y�s�Ӛ��䐑K-M��[ʤ���
�l��4��H��h��m�G����ݐ�Jp\ٹp	b8�_S}y�yWq�@�Hzp��;>�w�8}���+�O� !�DiM�J��*ʈ�.r� �Me���N�_�P��Pyo� �Z��e���C�����x�U�M^V��:Gj��u����;?��}��c�����C�v��'|~%�R^��u��
��<��R�"0��⬝G�!��H�xf/���'��v�*B�9�(�MHȖ%�ڝ��ɱ�w���94����p�, {�&z9I_���γ�ju�E���n�� L��ƗG@���+:t��5�?>빑���7+*uat��]4Y�(;�W�G�k��b1����֨3��&�	�@6^A?����hC��[�c�v�ٔ���3�E��"b���5;��He\ކA`t�ԙ~�ʳg �x@��PP ��>��'���R�k4�׆��M���X���L��X���4��B0\l�1����.B��nU�R%6�<��{��ߢ�r�
�
������kl���ҙ������߸� ��/�/���G����������(�u���Gؽ�:|�xIw4�rA�-�-�yh����aqg�(���#�X�z���/�����")z{�i����tuݍ;��MV�u�G=�Gw��j������d{�3&�Hs�NK�Yg�˷L+!�N(U7������AA��
?/�S6
�8Z�(=�n�6�r��7�|�����N���=�ӫzD+F�ҵ��Eu��S.��_�F�����mV,�2�tG���{DNU�ue�-��y
�A �?�a#W���擸�uFQ�uϞ���k'.�vg�)Pb/옫��:��?ˏI���D6�x(�|�8P�sK���e�榅��3ŵ�o��6�@�,p�)|�f�+�H�m]��n��I����0�+��qc��D�^�?���3�;�ia�]5�����-���j���U]�|���Y�� �����V����݄�xl�$n���gif�ͣQ�����'��mU��w �� �%`���Q����S�ec$��fH2�F���4o`�R��N�[�P�b\�/[�� \���� ��[�c�Zb9�b�4��S�`�t�$hm ��v�9�T�pډ��*��D���I-��Wz���H������E�����X�a߀jue$��x�7�t���fϴ2�N⛷
��]�Ei��)�� �~��'�/�p|A�
�O��O��!�s���B�����(6�R-[�9P�<V�Ռ�,�Es�ig��{𳃘�
՚���6�M�y��_������+�k.�8[�񍹽a��ۖx���D�'W�c1q�='6��D�l�4�p��OcB!͑K�3OnC�L��3�_�u�= � 4��Y���Ş_�����w->s]]=#>1�g/���>޴���<+j�ą�T��g@Q����I#�Q�y�?]��\�m<CYHL��2�W��l�����9�g�n,�D@{'BaPr��d�0�Q��D� N�b��)� ,:�
���.��TB٤L󓩗"Xy'9g�<ݗN��'��ޮ5���sf"����z*t�Ӛ��LG�/P�tmߍ]��cK�Z�o'՘2�I�� �S���x��IS�Gh��>���߭�,4%��x�6�7�z�
��h
:>�6B<A�'�5{�~5c����uDd�2�J����n܆	�N��hC'��vw��[��%�����<'����Q:��|�9`v�_�m(�
�
���X�o�[����� ���Z�����Y˺
~�fKg�p�7K�r����"Fx.0�_��2�M#�9���Y�f3媫���ݕ'�>��
Y��K���G4�'���'λ���V"��̰`�$�Ynr �$k�3&C"�2���}��U�C����f��i�#$�'%�z��w0������a2m'Q�[��6�W�ڽ�MYM�B?�\�gѯ�U���M��b̲X}*u��A�߉m�(b�)�
�9Kotm�?�z��V@�e�H8.�_Y0N��ЎR�A�jy�i��Q#��r��l3�_vvm6�2B����,��[�/�G���u5��� ��m�Ȕ�$�v9i�����͚�Sޔ�@��k�N���$����J�#���'Kq�9|)v_��^�����c��q�v6�c���G:qh���F��^��S*�AW�2�g���\���Maz��F���[Pڸ}�+8m6�Ms}�3][ᚄ�۾�DC�.F�[���+����d�}8}i� ғ��x��0�+`�W	�P#�������l��5�#�4S���ib]���%��5[cY��(V�e����t9�2&��0tp�Јd��|i�M�ò~L�q���[D7��S��9�����Z�b�b���2��V*�?ix��ꎆ�~;�?��os�>�;,����ܬ�1y�[r*��lĚ73��õF/��Bm����.W�߼���D}�Yg7TQI_�����)�ơ/ �V���߳�i�H�n)?*��b]!8�||�W�a?�vjR�?���),��Aږ<��f`���\�%��t�=Ⱥ-"�����@S��'Yjl�?���Z�hY����B��3�$��T� �@ tq�3��G�!�e�1�sʇ�80�A~7(9�p����`n�r�C)��	�?��{����YNOOe���bK�����Fg�w��x��罸��1勵zO$A��0�������#�xF�X����A�9�}�� ���M5�%!����d���dV��4�WW!��[Ī5.M��$��L�����⃊�?U^���w�c7�Ǵ��22������*"A�H��������0�Tο���=r�"����,(��q{Ŭn`��}�b>1��?7	Y�f�%�r�]	>2㆝3��z����-��A"��TQ0ԅ�	I&_i�d�}��+	�v��LdQT�Im4ؔ�-��rߎ��2����L�&�D0nDW���zQ�*�E��ꪨ5�,��x�xHx�<vC0d��B�������p[oO��viLÊz�K^�>҂iJ��=gSKKl���������o��V�&��A���2�Ί`���7~�&�D�����B)��.��'���N�<t�O�̔�:��q;���j��� �H<�Mk�
�(�I����;�P\׻�"�����c4� �)�)�[}��v)%�pҪ*��8�G���9�(8����=!�K �m(e`�Uq��Vo�J*f5�X1D��/�i>t��$���:��˿?��s��I�{ι닄9����ڳ�H<2'����>O�{ZH��M���NxH͊,��2��S��%n�vm8a��i�p&�K��3�D=̠RI�I͎�x�~���v Ej"�����#O��|�z`��Q�D��_���8	�q4/���T(+����V_���m1ں�#3TB䚞'Q:3T�t�M)e3Z(.�J�|lG�f��������7���P�ţZf|FI�y;��J쇧�s�|c��J7�˯�(+�=�����P�S	Q�]IΓ��i�!C�VhK�&u�����{ӛ�{��e��]xS�FJ�C�t$�7P���C��}��;�FLV��Z������7����ruPG	o��1?�R�NB��3��f����O��0cKбEg��#`ɭ�6�`b!)�4����;�fs��l��u2����"pwǋBU^�U�.�է��%5�����.js��/�C�ճm��)��/Q�����#�c��T���_�2m�����$��H&�]�pc4I�X�Zg Ƨʆ'}F�%���~�%�W����M��ǟ��j�L��Ő�� Ls=&���P��tm'f�Ey������^� �*��Ħ6�7�q`��웣>ʹӏ;��AL�ɻ{W,p�?����%:�V��S�ǜ�aº�.�_3-$�m��E��˧�U�6�	Acp���g�n��) ���	_�����ƾ�B��i�$������?l���9CmZ���ɦ)UÃ��K��e��#~�s�mdx���#6p��F�P��� ���:2����_��͞���*�͟u�K���5]������2��%@�nU�Db����|j��oӸ��b&�}����hr�ܪ�=�F�C�'=�Y�O��u��m첔/�R��3=�z��R?r��԰1U&����q )O��o��M?�$+�`P��drg��f�Q�m��,�X(�.+�p�<�G1^�
T��� @����p��!�KP�D]�fK��렷���>7B��C���,�|q������YGU-)���{�[�^2M��h�#	�>�"�'�'�%�e�6�k�iA�KU��P}`dܧ"�[D������J��(���M�DI���iߒtC��\̦2�:��u�eyx� �(i�dM�6�� 0��M�ّy�`F9hvmf�Z�I��N|����c|&��F���-u^lf�r&��Nʵ�^���X��6��~��;Z�@C�^%k�W�~_?*��:#���*����$��U׽z�p~� �b['.^~ D��K����}����GW��|F_a&��,�ol������K����y������B����Q�M���t�o����U܀f�Q�����SQ >p|��U���4�"��a������)E'��}�ܺ8��X)��wܼE��w�~�'��ޖI�T�NA>��F�k%܋*1SE�d?g�o*?m����愐���"�c�<��SLyK[ �rN�}�I`+����P���q�#uv'�ƙ^0�}3�� gU�Ů�,0��cw[��J���-ْŃ��(���ӈC���	b'b�BlN�;#�ۚ�64g(��$b��,Q}L���t	��і�8Re�wH�I{q�=��u]��p�fB�@Vc�9��W+�� |\�SQ�'b*[p��k� 5�9�U��+{���^��[Q�q��۠ gcF�r��-��q�O�3�_���h�ux҅��n�,��%���������	��r.1<�=�%��|j9�ǘ��h��N ��C��Ti,��L9ij�J�J	1�׺%:��O_�=+�U��wX�?C�>[S���3;u2)���>�4�e���h�}�Τ=^�T���gپb��m�ؔ_��쭫/�����*�#p܃��)���?��QC������=�̳��uI����A�I%N�d�W��s%U>^m�U�N��q����r�?C6�cV�G|���?�����3���l�B�J,ެl(��Vt��V�r�vh�59J񄭞C���0o�V�"�`�`7�i�� ���1�����SZ���V�Qǅ�NQ�((MW�k*�˂ΏS��I�Ϩ�%~R����v�������";`�4�dp�Ȥ(T��[�(��19B�>��#U"�Y�s�x��`�:#���,Ь�سZ{�_�.iLY"�j�o�?���=v o$������ y�8�:0�t`ò�Y�$%�R��I��!$U��l?��,O�4�P����|�o(ɂ1�,sN�*�����L��D�ڃ��d�[���>Ԡ�5o��S��j��΀l_C��F��I0��L��*,�t7W��]���q�����(�Ja3�����I��_�u8����q�5�~u2F׺��R=8Q�w���5�;
�س&����A$��d3<G� ��D���sc�����e	�Ԃ��%*��el��"���h����xG)/*>���Q}N���k�*���7\}ie]���g��M��`��9��(N�8Ҧ=��X�٤���X���[D|ᖨ�!���ļ�E`�`��R>��:��������I��&�p�Idȉ�
��6'M[���yr[1��N��C<K���w ����7T$��1��e�=�����f��Mc���rR}Oju�N<���qL8�`�H|1�<��AT����Nn�h�K1f�_5�f*���`�Y508>�N_�!Y��'s⥌*������|rRg��m��+�3@G����Z���5��)�G4S^�}<�ƍlw6�+�u�\�T��\x�F�"V�����I�_~b/�.���=�F�/�\9��̂c���$}z���{�o��%�V1�����֭cS:f��������I�x+�4������0������7	t��ey��se�hfj7g�Qa4�**�)���]�:U��x��B�}gj� �;���*��s(��ʨ{XD��mIV��S�:'2m6/=�%�}��ȐҦ���]ȫ!$1�ZT�a_�
;�(N��y�ݾQK�ۓ��O��# f����>!,�;��Q{J�[U_�.�w�y����9ơ�����S�.l���U6��t�>�������^Z	��Z� 	�WՋ�l�3�_��\�uIX�
�?��*J��G�M�1���7S�����Ҕ�T���ʇxk�g^��P���V��;�m��s��� t��52b�z3΂���
P
�Ӏ26��BU��  (����s�Y�]�P�x΅�^�J�"���e�1�@���H��U�����p���9e=l�C���������o�y����5���4W��͕t%V��	Vr��Μ��p@�H�c7�g۪�z�ґ��|�\pj�����d��$�`�9&4��Z�d�rZ�]��
CN�zI��+�n��"���QXM6�/ș�br8d�*���c��6�O����M���Ǒ�������)�{́�7r��Ym�'qF�={�G�7%�L�YjR�T��q%n��ù�gU�S��?��u�����5���1�`�{y�)�x�0B�� Д�I�~�~L�P�'��͞�y;&b+�$1���N�
đ�@O�E~q��!{g�I╜3���\����"�ء�f�l�J�*<��*4�fr�O�z�d/�nu�tu~�(':9yV�_,h�� ��ȱ.��L1�ƿ�m�3.=����m4�����*���Q0��tsR1�9�X<^��ֿ]�i�5��ϷA!��'h�%�R�Wr5W�聂�+<�!��O�J��M�(h 9ote?,_5�"��2#~�Y�X@�����ת�o��3 �lGgε��eV���ȝ-#��hu��0^��X�?q��=��}'A2F`�Ǝ�W�����IG�-�<��;_���_��/-�	����o5��z=�T����2L���TY� E�i��a	�AD&T����*�ы��9����J�׌�.�ʹ��`fs���+3�WBM:���-�#�?��u��ۣq��1��.`�\�⛆Fğ���y@�ؾ�����;%��f�s�-��!���F(�����Aֹ�z���|Ҏ�)��;ji���k\��������Dȩ2ۈ�@�\�
7��/g#�F���&1�"���o���[�2��)�(��K�|��귾�;�.��)�;�zOA�[���S�?d���kY�iO?�Iv�irL��a5P����/Ȃ@��E�$�4�4zf�3E����;�VsA��lDә�A�Kp���:d�J|)��s���}G�eB#k��_!:�|G�(�UG��*:�CS��I���KK�d�	���B d�i�'�7 �E[�]�����'�ά��*����e���k\��t�'�/5O�����h<E�}�&Z:���q�ë=���.����~뫘i��D�����Ҕ��q�U�*P�����pc\�5|����#&��[ٳ��t�⠢��S�6	!8�^+�So$Ɖ9IG�	�AE�[�T �^�K}m�|��F��M�^\��O��g��-�����VU<5�0� ��{�`]��J]��PW���$���̸�}Gk'�ݎ7�j֥v��$za<��J,8��1-���xx�	����y�A�ć�d:���q>!m���/� ��%\���ev�\�ڂw-����Q��S��5���_�����)نrE�r�:�6Զ�T�Dٝ��h�;�ndN��"WI�o8�L���\-5�s�գ���\#��`C���s��}K�ͯ2�Ae�)W�I�d
y�,薶�Ct���s������7j����Ua?[+mE�ǫ�����]�u�a��;n�M@R����ɹ���>Z��+8Sm�D�2�]e����+W�6]��+�L���z��B�o�ׅA4���뭰�oBR�V�YS,�ϑ�	#Ve�6} �]t��:5�j���{�_��5����h�&Q_�]��M���
�f�ę��YJ:�]��}��+%�Fj~W��>Kz$.'���9u� $��
��"V�w�[�Qj���w���<�3=�wh�iI�Z�o���Ž���8N�" �\��s8ۂ��|�v�u�3�5M�yߨ��䴧ॲ�x�[���7�V��T��.47Aq�b8Dw��e$���{L�g+HE�S0I�o��4L�H�r�s��}��k��=c��>�O�>q}�9�3Z+F����-��I��B}�A��]���{	Ɋ��:��-�Ewݱ���:�N2P��Iֱd��ɭ��]�(�ߡ��鳛���g��~�&eiV�Ox���V�qƆ��E=�j�����JF��ܗb��� �;��DeM,p��ZnO_qA��LV�����9Fh+�J�(�ll �R2y����u1䶕�%�F[�U���݂����W�K�(}�?w�
"F�W4Jyg�7�\�b���b/	o�V)�Mˇ�'�+�v_D��Zh�p�$�L���}6L ���ֳ����ꓑ�-I���.�r�V��Z���ޱ��5۴��6]e)M-|�¿��^�����/�ۈ��Rӱ����2y�����T�s�J~����^���� ]jg�ֺ�/w�֪
��N��3!k����'Y��$m�g�)�RHE-���s4)��~� ��Pñ�p����i0�t��G����Vhp�}�z\�s�jo���Y��2KvW6�Y����-�R|�o�n�6��a�pu�z"�m(+@��rS����G��qÒ�a5-����M��	� _��N����v�ζ��*g�����܃s��;�g]rW���G� ��D���s�ȰL%ǥ�&̜�����7�5� ��ϊ��И;��ɩf�4�R��@�A�ҞI�GH�P���{_�[�ⷴ��e�!W�_�	<�>��*p�oX�s�vO}�7
[��;ç�h��4�j8�b��;}�o�efC�ŵ�z^�ؖ��j���۾����9�x⩷���E:ۺf;12Q!|:�?�G��(+��<{�Ք��K��֥��^����}�n�\muYH�^֎�
g����z	�U����Q0�(+��|����qiy�&�m������J�� 3�=��:�,�5֜��f[�ػ�1��0�:�n�E�yi��������t� L�5��0�Yk�z�1��_D�Q���Φ�:���u #�Y/��_�'��܌�G�=��.�g���~e7������%̈́�)̙�l��%I�?@{c�� n��L"�4г��Ơ*4Tz@�P��i��8=� (r¼,,�+k��7�Gl����%n�H�x��e$���nAs�h��#����c\V|�a�JTi��!��C�ߢ��H��&��*ͪ\;�9}Oq�
v�~Ѡ�܉+1)J������J��]j���=�c�.��L�4��)���%U��.
(d�� ���3��'r�	��L����d���Y�E�t���7�_�[��M	%�,�`ʎ�_����wxڧv@���^:=�������ƀ��ͨ�xQk�q�m���,�D\����y��$�F�᧣��mM�E��W'Gڠ)H~���
)^j���$��Fd4f��I5�� �����!;m+�m��85#K���f�s�/���#]r�ɻ3��o���V�}/�E�c �4N��U����1 i���ߨ�����;�G~���̮�X�'�<�ۗ�g�k�Ol@%=�Ƨ.6��#m��$� ��°KEZrOzlp�ݻ��{Q ���f�(��b�䏎��vm�ȍ �\{#����+��S��X_ކtL,c��(4]����`��~�N�k(��<g� ���*CGPԇoX�k���5�� ��W����� �*z^��=����sD������4�BU�t���u�a"��	���Z;��D&T�TJnB�i��>h����S���q���(��V*:}��S����@./`d�?�Q��o����h�+'����:+�1��i*�|M�HAO�Lb����w �@d�JV�.�y���d�9���nF-ܑ�ʏ�=S�a���#�9^��j�D�@��f(�"ǶUJ��F�E]X'cn&��ڟB�#$�k���TK庘��R�;�s0l�ʢ��ԨGI`;������e!��9���(i���d�&*'�z��#�J>s��6}���lD����:KE�x���-�@)��ҥ#�M9$^����ٰ��4����g9uX��y���|� �����9d��H]�-zS��F�d��(BpJ�+R�?����$4����g4h`��0�2�;1��q�� i+�h���p���\r��S�ҿ���<��f�U��i�#�
���M�S���x=A�����_>
����)P��h��(��}C�b��69��l)z��#r5^!r� ��m�_-�z��ZV��~�Fǖ��5�3�?���۫id��
eh4��'qA���t�W�VG�z���af�.�	���V��j����~�z��-��I^B���t�b��zx�?O�pq�Myh$�5�i��u�׸�|	������e��Rq_u<�es���`��I��%����f?&5����E:xcy9�_2���T�[#@T�c�)¤������%Y�� ;�h���PF\r�؉�0)`uޚ��� ��&@
)iE`�#b����]ET1G�T.N�Y&)�߇��W��B��Z)+�
s,<�is�u���HQ�<��vQ(ʿW�\��Ң�6L�n����8IP{�Ыk���������	��d��z�t�AO�Q��3J��te!N@FXez�\�l�wPL�Q2?��\��1�P�����>��?X�2=��
v�8kH�@�NEG��ѱ����	d�|���$�)v}���CC�9rN�ߞVXdcsw�9�S�ss�Ll�{���N�5N�k&�c.U��|f�2z�m�[��0e.� ^�Ay:w}w�dn���3�v%i1���;W����Q+�W�ʜ>�hSo���f��6��^����]����;0x-���+�����Ҋ[�3_ V��x� ϒ~j����ψD���M[�S �ّT�U9��(HU��$C.�C`+��3��6�)�F r�.<J���x��	�,�dP�%�� ދ�{�3#�N~�%
�)���n<j6nU���)��ݣ�]0=��j�X��
v��W�"(7st����@�ݮbƑ�9��ۄ��v^��M[���-��"�
d���O�����L�i(���]vѡ�:S,��D4�ă���2�Ch��&RW�I�KCN"����k�Bz�����Y"��|^v)�@i��z^�!"���u��>�i� 7l����U�3�Ҵzů�2��I�uϒ��Z/�I������������H GXî~�Zn�4����kt7�	*B)�����I�@�\B�2���t����I9��9_����^O��S�\pV��>�(BL���m�W���������XSJ�y^�CC.�%b�*����5�ZHv��{��U��37�q�}�cU�-���6��HR���.�6YVqj�ܐ�Q?��[�5�֝Զ[���I�Kx���wM1��#O�ua�� ���Z��e��k�i�-P��Z.�����w�7<q��"��h몦�X�;;gkp��&V�7fe��V����:r�X�~��2�}�@J��[���z�(�EՓ�d��p�a�=���Tb}5]u�[+J<�p{B��-Uw*�AJ�G��6.v,ȏeI,1���$��]��`��3P�J�K#Lm��0�^��(�|.1A�;̮��"y�eA1M�{M���@��aCjxq@g�d;Q�u�Q��'_Q�V�r��<�uG��_:�:L�۾�Kk�w� 2�<ܰ�fK`Č��Y8��\*Wa���)����S�_�F�J�C1���"�r��� ]�_9��*f��A�J���y�`G�>h�����I<�q�<$�D4�3~=�-�-5ɤl��mr�/��s=jο6��1�dA�vמ��%K�8K��vFƂ�!�#=��!	��<�G�z��ý��埩��(,�(����"���un���E�{~v�NA��3S���Ƭ*n��� �y*��_v�^ò:Y~D����َ�5�K�U�7fZ{����S�� ��������@gQ�2���I�g4��g9���ib@r:=�� kʷ�z?̓��0��F� 1c��_�
H�v*P��9���Z��du�J�F�1U�	�MZ��e�!���Z.��ay�k��c8�čj���FҢ��ls4�d��2l�Ǣ(lC�c#���:c��V����7��9$]�gFD��D��X� z��<"e����Ǘ��OD�=��.X��bq�dqҷ;+x�����;3S�������m9,Z��qP��=���l�a~�s�uP"�����h�h@���j�ѡg�6U������.�t3\������m��2�=�0R4�
ӪְV���$�ĸ|���;�}��dYxs��o��A���6�6#.y]ā[��M!t�1���) �Hz��]w-�:��m���g�A���$b��X��5L�sP�QqB��s!�<rW%�g�N }">�7�O����yG�ZCo	E{�[\�w#�P��n9�#ҩ&aШk�~�wֆ=�7~�EG,U���r��Nnb@7�yw_���`g��,|%� �j��z]lF*V�8lI�2�2Y"�,�ً�c�eF> ����	C}X�<�^�׮g�i }��(}�}�8z�g��_��-�l���+v(nE��*d��e8^�zA��e~����R�A�&,~x	6�w-�B�,�z��W������#)T<D��x��j����)O1�X��:g���-�`>��>��x	p�%��l�u�H��E]��.�)a &��� ����3U�IgIf��D@� ���.Wx� �mIXt��KU �ě(��(&7;����eO��� A�������*@��9������ƨ�T�G"$��1i����|)�JM�;b�ԛ�J5LБŀS��(Zt�����tǟ<�Z!� �0H�/�;jc:���p;]lsc�oͷ��l��#L�CP+�2��%��>��z���rGX���k�����
�hڱ�� /���Ůb֋�$�p'@����	�wP-�q0A���`I�T`�ۺ��@���.��~ �ŢO�_��S�ȩ)=|�T����=�����?ݭ#������W9i^�}0ƻ�*���2����p&�}|E�Q����.�*����="{40�2Ĵ��E�T�)y���1�;(I�/���{�Gw~��l��('���:��N�S�� �v���_�����O�Um1�g{�:��R�-���:��+�0�yw�ۂi%q�m$�ن�ԲmĽY�]\\n"�'��0f�Z�{%��\<�3� ��L�]���#�ݥ�,��ř�W�f��,�Ö�~g��)�׆Nc��PJ�J[��������J� c0r��9��O��g���;t����ƥ�����¦Dj'��J�ɯ)��� P:��}��c��lo5E���;���ӌÑ�4&^S:����9M�[�'�F�d8K"$wbC�]Ǣ1�KǴ�,F�$� w�ҢbP~��r��s�X���$���R5s��*���{�7W���=�˗f��;\v����zv+gȟP�{��/��im2E�qc��ŵߣ�p W��$�� ;�n�D�_�դ�B��[2�±�M����7��ݿ
'�5�D��.PC�����^��ge{�>*�y�<�����#;䲽�"��?1�F���8�?x�I�-�9�3w<"D�a�z�?�>�g[\d���"���	!��Ѿ�5h�D?�����,���&��&+�|[����J�b����`��0i��m�~��	�ê�>�x�ۏ���Nh[�����b9ܺ�P�|F(@�>M�Y.�"��q�o��Ȗ�;�zD�,����'w�R+܊��Af��>͡p̐m�>��a����h�������S�Ǒ�ԋG�A^���s���ߔ�_-�u����;&ߵ��0fe����s��:�7՛�ޕ|@�m�I���0J�k�A�d��	�ρ����9�	�"�)�\�kwfՉ@�p�'#��:��#���:��a�.C��u�D.�1$���U��)�w��m���;@:����� �vq4����3��(dS�pH_�x�gP�ǿ~�(}F3KV��e� �}P��FƐU�"�)O5�?�$��5���7����_%�}�]$��n�T3c;S�Ӽl�-_DLL�dzAp�~��閘�_�(+�)�Q� �y	�$�-��ے�h�ndԖC������$�C��2�F�%�Y�'��$�3�|���C �$R���[,�Nj����8�v�����6�|�~}N�.3��`(Zqr�ݏ%��u� sx� �ϒT�T�ܛ$�q���0z�>G�Jˍ���~C��_����?
	�+��F�K�<�� ��`�d���2n[�7�s�]���U�,�k!���0ng�^�޷Nqș���Lw�l�ob���e~�����L�gAjӒ��#:�h�z�|���p��(�eQ?NG�����I�(�p A�6���SUB���[����p�A��䛮/?f��I%ŗ�v��v+<L{'<*e-����j�������/���7H�:�Es�Q��!=?̜e�
U��m?��T$sM�rM�5g;�f�<0��>t'�3�;&����6��?NP��d\E5�\@)�_ç��S�8���x^���Ds�~�cҰ Cpz��z7���c���{=�\��cŲ�,���6�3�a �7�IC��6���V� 4��*�z*�;�v��k��3u{19��,�#����-:�:H�5�v4o������q�]�y���Ű��o�	���
���Er�4���Ad��É�g�$sǽk�=�'�j��s.]$�=��3��$�3c,k���V		��u��O|i!Uy�]�F�aG�{�Q� ���9��;�T��.�>H��}�N8ޕ��#&��˭4��C���r K�si<��S�#@Y�=����pt`�a0Z}7Lu�aRB�=>C[��4�3������hYց�V�-�ZC����U�l� r��b�N}���p�đ���{:-��N�۴̶��8��ك#����<�9�'��C ��9��$�c�cׄ�^�JQ�TddWk�΅�FDW�$��9�4�I��.?]��E��z}H�E�@v�׉PC}t0�Zb!�^�LB7nz>I	�֏&ƌoCU^f�H0D��.3�K�!|�{��(��٩d3w2�JB��BV��ZE�"�ܧ����S���PU�R��d�F�5�_x��L�?9�SX̷�Y`��3ܡ`1h��IՖ�Tk�&���K~1�.���Zi�c�`e�Da	��,�|J��x��ƚg*Vu$Nn���97��@o�vB��6�<�xN��W�ߡO/4�]��	���b�9�����G�=�PUa^q`�i���]���~�{�H�B� �6V����xmg@��'�ѷ�޷K��r�i7%�|%Jbl��
�`������Sڮ=��
�>�}1���(���I�UeV�b�	x?f����2�xх��+��ަ0���G���ק�|�ɥ�T0��7&�2Y��Rk|�~�8�����bR��T��f�b��ov��bcz�\
��3���B�D�V�2�F}{-�W@�=�0~=�M��<1=��K� �(?�a��W83�$�,��卧i<7�ba#�?J�<����B����.����1��K�R�!k=c{��>3]O<߳P�a��W��S�.�����ut �V3�ⱼ��ǳ�m.V���sH@�vtq��`Uȓ�y���k�#��\�B)�Œ1L`�5�3b���Y��i��f�l4H���Y�#9|j��)��D��\�1�8����&��D�Ҵ�^_�����Ѧ���L�b�]4��N�*��y�G�@�xn��X���8b*� n�����h��1�4ߓ�����*p�w&V�U5�=ʮ�
5x�o��$EG�~��n��6V;)��#<��-I{W`P{�:`�C�	X�*��Աc�V3Y�<�Jp��
rg�܃�`�-�P�Z[Յg!HS��Ԛ%*��2�(�$C�kQ���"��~���v����&8��ʞ>	!��3?G�2�^8g�l�F�_d>��53���e̝b��O-P��'Na9�3|�~���ؔ���T�\H=���>n����>8�W�}k��?1�4\�HL���Wn�%Isq�xWe
�� �`��a�J�`��QҼ�s�%"� �CB����h�2N�3�j��~���1k�� �F�bê)��n��������Zc���&�n�Mp���t��3��h
�f�5�Ÿ�
&�ג�?3��=������	�Y�o~(�^[��\��kZj�/��;�Dk��2�J��E�"R禹}���8������<����1�[h�;Fp �҉^�SR�K�Jh:��m[Y#�`�\��cV�-�P�N�M��(%�^������S��^-YT����<���'2TV�f���V�,�9F��J���o��C�"
Sy�S�x�+C�#��UO�7��n�[�iwe�	28/�o����c��}⌸�V������@J2gT�
pC��](<H1�����~�em�D����؎�ݠL[��������G/"�u���IZs)�3�aˀ��G�D����@�^�i���jS�or�(
�o㩨J�&|���ή�n����fÑ#l\�`9���s�	���F7�PA���Q�Oh������/�c���:����Gϙ%����$:v:T5zՉ��]�q,߂rh֡<�u6�jN�i��Ѣ*�N��٪dW���=V4�pڼp]{�����Ⱦ��<s���B[���z�+ZŢ��.vU����L�{AHW�'�%��g'n�δ��Ua�X��k�ڎ	(���=Բ*�=��'Ck"4�?�|��[���������b���X��i�J��£��� ���`O���m/�*���#���A�E�Hb_ᆾ���I9�mDR��n@���M�<Cj�e�\��/��ϵEwA�<D.NFLUXxc�ǲ�E����
�g����F�!�0=�� ���Q�ϛ��<?�la�J"<Q}P)�	�SI��)0ǣ�������tMI��|Z54����:���Q�����+��4��J������f==\؍r����uo���y���� Gt��;�f�|�����u��n�:&QBj�9�ht���#е����p>B�LOs>Ό�nF�����|���f!�*	s�"��9����wXT��|�|0P�0o�ů���]Yօ$
�
"ݙ�{�c�l�P�g�$y~k.�H��t�C�#�pho�
�;��v�c��[�������+�%x1V7J��l����^��$:�g����[��Ķ��燹i|�b�����v����.y���LM�S9��^��KM ��@���{�����5�;��U�#����(�{�y�*�j��{�G�*9�����G����W9�ufO\����G`,.iW�}I?��[�`',W<O�`�6�Fg�_|]����u0�鯇���ӡ@�y�ڵ�Q��ڿ���@V액���MYx|�y���ؤb$^`������ը�CE8��� A�+U)��\��y�6���
���A��U?_�2�"���<���1V?Դ���V�ʑp���@�+oQ�ȕ&�n��P������#T��|OJ�*����v 95�e�����	�}����[h�����๒�T�qٽ�&	m&Mҵ��QnԪWޱ�?/�˳�84���UG*b�o�
����Sx!�	R���3G!7�V�h;��?��,��^�H��/�/Ν�9�f�`�����+p,mu;|�SOg~-�3�:�"I�m��3�j,-Ԃ�-"�n7�(���P6Y�]b�x�Ay=L�p�C��2�;$n(9�rMHVG�����;�O/�<'������eV<�"հ�s����H���Fg� 7r��˄2�S{�	��.��AF���+G=i�G�J>����،�fCn���#�#I��ǔ��]mR0S����iQ~ѷ�S7�}Ծ�ԕܵʭnm��5�Bǉv�k-*2�c�>ԮB��o��K��@��n�;d���XW��Ч�YI�0���E����_�d00fӿ|�Q��:�����]F]R���0x�-H�4و��}t�S�QL(�kP�9C	���hM�_'���9�$��^��$|B�M#�Q��HS!-}t�Zh~%/���Rn�G�L�!5OH����|~�՗S�tՋ�Z����0��&o��E��G��\�;���I���+؄��L:2�Z�S�#���2�_4�Lv$���x'v�݋�M�^�ʈT]*h�֖��zêF��p����[�u�h����]U�XL�E�|���Za���/��]�3�^��p�C�4�E�?+=�E�0����y����������RT#�<kS�t�Q�U|��6֮�m�ѭ�1�n�-��U6�_�Z�h��0���=�Wg��.���XQ�����=�J�T3�y���\j=;^fhf�{��5oB�al7�8F�-���8���vדZ���S+�r�I�n��G�gN�����)L@�(􀲸52�u�@�aBh���M
�j$gk����ڳ&�]�ZI7b/��K>����Ru�	�z~��7>� )�������p�&3�9���y��\�B���Q�-W!��k�057_mT�]�>��Kһ��(���Q1��wm�疦��_�6��n��u�ޘ��Ed��u��R����''��R�9��s���1����v>�@��Q��"Z���I`l�(!�ʀow#I�g%���	�>�Z��Hh�L�m[�7���Q�E֩:��sD7�0�C�:��JR=UIQ� �K/°���:�-A賿@>>�-Kl�ǀ���:�u%�	�7������4�7��n?�Oq�l�Ud*{�U0���p
H8o��:���y)�͇t�?DZ��8�h���.d��E��NnRFݴ�H� ��?R5�a�~��q�k��GU���K���H�k2UE)��aOm؋V������[ߖLP�W�C���^6UܹW���x��S�����8�wT��m ��K�gG�
0����, G"�A�j���j�"y�sx�'i$S��ZY�(���g>�S�f��%�[���a7U1���5%.�n�i2�XH�%�I��C�9'FB��r�$?��	i'��Q*�T�P�'�Zo���/=�����B��z˴7�~��t�+�%	�zb���3͐�0�wc4�;a�1'��of'��x�Ä�H�X�+��I��h�7|�4�(�8\Mj�E���O�XL��E~�1m�H�8��tT�C�t��'2��ԥ���(��x����;��fH�����a���XPɸ�M�R��	�G�����Zo���l��oh�ג!ֿ#_;�Ǝ�I�-�I���mf?BV>�qP��[߀�������"o�~��:�m"W�I��oQ�Q�shx�����Y�Z}M ���4��=	��<�����z\�·w{g��hH�����ǵ�Ʋ�P���ܷUM*gH�!�4ӑ/gbG�7�5`��%��Īo�&ܿB����T`婒V�g�`}�0ƕ!����csY�f���Z,�]~`�Lo���D���-\>�f�L1�jct1����  �~�w[8`��DW��A��e~])��|��'p:�M���^�˞&{�`���5^����*(	�
Q���<��C��m�=l�/�F���p]����e�87��`6G���c<�������p�|��?G�mt�l��f�#�����'R�=��r�>��4*E��]όk0/d�s^�2�Se�Ly�]��Z�e}�9]�Xx~+�f#�C��s�-kۿ�=S���,�8u�<� ��c��I���c�K��1ңm^�u-Q�*�,E(��hp	K9V��̸�M�֡ĸ)���*g���3�f�L ������?�h��6���1�x��*&��ƞz�5�D&��;����z��,	;�c�mV�,0?]�\^�h��뎀&����"W��@S��bn�k(�ܗ*��CZ^6��îO	�X&[���'�,H��m�<F���a� 5s
X�p��
b��񃐂X�ZN�y��AǈÖ����f����wNl���󸽸�C̲ɚ��BAʦ
��3r��6x�:�u���h}.@"_mt�DT��IŚ���m�蛈:���/9�r�_(���D)�݋�UR����T�x 8��e�ZT����C"��:�*�e{�	���f��?.��v��pf jB��Q�2X��}�Z��F���� ~&��_��^�+����0���AӦ�2F�I��g|�_[���P�#'e2W;������+�S,q �Xd��%��@��}��t=:VS7�
�/�`D`bu1P��W����8��I(�4��w�e�����*��U��f��1y���qHzf$<$D��g7�mW�2�"^�YU�ܒU�����H�v��P��|�Z��)��$j���fCA"hƪr�@�ʖ;%m�ڙ&��I_��_ �q!�8P����U(��S�NP��`
�ucy]�nl����B��`�k��ї���M�4�R���kX'��.�3���e:��R�p����XpLR�rT蘇���*���nLq��z���P�m�EX��X#�q�$�q��ۼK��j���$��XQ�9+S�:�o����݉X��*na�k��q�'B��?����F����ݥ�RU
�(o3'���5ʑh�<!`����T��V9K�E_a�/҈%�@�q��nF��]�h���_�ޑ�~�e�0�-�YQ��>�HZYe�E'[��i��{�4έ�<Y�ĉ$0����x3F��W�?�>���s���6�b�4��꭬���Fl�p����ux�4�Y&�>br������z�H��reˮ�j�l�H�&�F�A�����H�2��+f!�$�L�G!��z��;�.���N�p[O�����$�|��@����u�%}�*���Rm2�N_h�F,�,�O��-��������Z��/y̬R��#�)���.��܂ȓI�(�[9��)k'�5v���j�с�$��we��<m7Pr�	�A�4 (CJ���00��*�l�|��e�V�;[=G��w����9oM �}��Ҵ�k�<���^��ϯ��ֳ�Sq��Vl�u��+#�*?�\>j�����[̅e&�9�U�9�v�C���1���1�A<?��\�7�^[t~�U���7��ڙQ�٪L��kk�����X*T�ͪ/Q�	�l�B��y��]Fg������ ���C����g���uG�N-��q��/N��;gam���`�(G*nl�n��5A�wo}���X��3�~�t�s�,y���+�W0���K>I7�O}��#�л��ܗp�p�&���KV�� 3�$�=�f~�{��4�S
�2��#J��?�i
�����@>�4:�Фr�����5�I(�\���d�E8HT=��o�!���N��de(��s��Ӗ.�	{�"7C,fZ���)�F(�r�#�{pF���q5��]�%M��;U�C;B> 5táb"�����7Z�����l8�g�LH���A� w/��� �+�d�/��s%�R;\��}(��EL]Ή(�e�Ք�����<���������JyR|�S��lLX��p���b�q�)�Ƌ�/��T��jk�9�aDr��r�c-Y�]�@�����J�o���p�DG/Bu�B2�R�~�(���?f�UC\x�V�� ��	��1��灖�Q��AAb��[C�<"S�m5�Pg�b����a6�:�7�*=�r�^ťK<�����H?~�:y+����x��ff����8C�_����C�g���+�a��ڲ�L�r�}8F?��_�����u�#�mN<o
hyRS�`C/;GMsZԬOHE!�(����ue��6c\&�,�I���`�Or�|����K�q��� �!�~Zu���7������a���OEK�>WY�d
�4Y�_N�udcĖ�뮄���Z{Q��������-98���,XrS�h\oD�q9cL�]���hh��33$@��vo���� �HP�M�k�yZ�U\� �{ϑ�S)���IR�����}"c�Y��)�˄�.���h���"��y�ZC�Z%k���?��^@�p[�2�i�� E|rg`�
� X�JY�$�]2����H�K��
�op��~�@-=�x����(6��y��u�7�������p���6!��dfg��t^�4�񭜗�x|y�]�Ei��'&w0�n/M��f���:��{�tO&�b���Xa��#:��0��%H_<�-�!��Z�a,��-��]p����t�b�i�l6O�0��̄qW�Gt�?R�������#c����qݚ���a�}hꧢ��9����˿�1���C�m硷�[�B���?H#e���^��o-�MV@��!��V2�me��@����_���|��FS�a$�����u��Wd�3�]c�W��Ă�Z�;��jp:="鮑qe�����N�V--G�p�OR�J����R�?&A����x�!˴(��
�ӻ����2�4�q��Q|ɵ{* ��q�K�#�/�Ni,�*?瀒J��g^���"I��@\K͵:��`~���8�e���sRږ�/���ؼ�r�
T�O+���jQ�7_9TG ��L������+O���z
�u�Z�%l���É*pN�X��'bN~��P-��:�M���{X�,�bq��x׾?M��~�YAF*+�2u��������D[�]���f�x��e��v�|�+x�d���#�K<�$��*\��D����iRoh0�XqP�����c�%V���_#�9��⋖i~s>d�����G�jJ��O����_%� ���H켧|�@��tb�n����؁��þ_y$��� �ؾ7'��O�� �(��3v���X[x�����Z(h�?�%��0,"�3�E�:Ўh���!K�x�t�l���?����C>Pķ.2�����5��jt�@�ʝ}��7F��2�� �<��,����ڹP<�PlӿH	�̘�
��~��>i���Ь0ޭo�{��Z4���:�s����h��R2�S&��hU� �{-�~k�E�$��ҝ��{�k`��[~W��E���(�����|�!-Jm���a�{���y��¦�$^[��wګ�IB��J�Gy�;͙P#��S��"��䡗؄ _tGB8�y)��3,��;�J��{k�=���]'�;��8��B��%���	ou�
gf��W��c��u�V�[t���O�RN�a�m���b��������q"�Ry>�7 �Q���Z������OU��dۛ���W�t��9c�<+�Bx�k��eчL����.)QC�o#��S\D�ü����.0���*�kU�C\��uu#W���:�n�G ��R�"��̹In�a���+e���U����#��3JOR�\K.�����U;5S̅����z�����B�\$@S��n�5�)��4,����^|�J$�@�z��nO�.y���%�~I�'X��`	��:%�<�3���0E�SO[�NطwK{<�Ȥg @J����_r�9��e�;^�����T����v2{PƟ]s;��v�;�>�_Q�3�XG���H���x��zf�� ���Yʽ�om���k1	��9���w���a^�H�#��֣����9���h',=��b��9�O�N���z����B=0�ɪi�7	��y��P�h�r3ح��d��N�08��4WŦ�1���'�I 0�hqXn3��ʢ��z��[�e���J�^��$uC���VB�����o#��L�lS�u<M,؟��G����ҝ����N#3��EZ�������<�S����k�uN��ž�~f�A�� �gG+]�K-��}j���l�3�]QU��
�$ר2~�_�Z'yu�U?=�c��?�S~��h�����@�E�|�0�b֭59�egv�ЯĢ�bT� �@$PY���B*�aυ	�+�Rě��p~K�m�mތ�i����� g��4ʆ�m�PR����{N)��n%����XɳC���q�8~��l�5�r�WAsI����sm���*�?�Q4�-�x߹!n�e�8�e��s	�#�X�
f@��B������W���L)�#�Q��xNTT�l<`M��)ҡ ��#��bE(��G����U��xDS���t؏�yl�%V2�>!�M�<Z��PowJ�y�4BSͽ�-�JD��E8}�Bt�9����í��ߴ�s�.1��Zť�^҅I�Ȩ��|��,�����n��Z�ဌ�����5���u˲����8�=˼����<�p+��P50�UT%��Ux��}��Of8�>g��9Y$	S#	��1���HE�e�/y?I�TsJ'�R�����&��r�O�P|W*�V �)A�c{`����!D�J '��{sB	�y����$��j�`CM�Jrwaf&�-H8�x@�Y������<����U_N;�0��͙nB�u\�w3a�Q��'^Is�gE`�T4�y�z(iV��7�/�>�y�W���ɔc[Wn�&'�NY������J�E����Q�g8\���뚫�AHM��O��X��zR��ؒwk"(�d";���X���Ra������<���{Tj3���?Ͱ߿BQIu�#L�d?�����I�����Gu_�1����'t�-P;��^����)�g�K�c�����ڮ��Ⱦ1 B/�5=T,�U^���0,a�G�A
._��3-�@t�XU�=2�\|��E�B�bA��vk�|�f�[�@�4)�#{�� �k=VL&̢��9�� �
a�[�;��A�1�*�z�!�΢�#�ЅK���җ�+���2��{���_#�(g����w("H��ѧ�5cp�߿��\�#-oF�r{�\j�	"� �1����6��1��2������:�a�ML�� �z"s8{��4��S:�ߐ�v7�w��%׋ u�ԻbVrG%|Ҕ-	b�d�?{�P�gF-n�z�L ��;�r����m:�:J����9c,ҏ����´'J��h��<�X#!�D�9�C��n@?F���q���1�n��K�{�6��*ԝ1P��J�|aJ�z�>Xa������|�*Q���iC�������I��ʹ�۽���N*���=y�m���7�n����I��کl�󸬱[���ب��[�D����2? �q7���9�c��*m�B_E<[�1 �;�HY�l���хP'H�ȳ]�~��\6��'���ZG�kb��sQoh���ʾ���G�O�l'	N����4�ʶ��37��ܯ� ��s[�A.�����?m��]�*~b���_M�:q�ʇ�pB}�<]p�TU���,�&:44e�r�o5eetP�{ν�jZ�8��ZY�OiE�m0�����Ym�M*���蜻�@����>�Q���f�L�.�̠�p����>�pJ+����>DI�i�EP����P���.H�Kt�4��{>Y���REJU�{j��#�E�J���>��IsA��l��_7��6`�e/��Z�n�B�D���Y.���N^Y�x�B��5�h(P�O�]�@K�Sq;����Rɍ?�|�m9<^�Zg���~Qb�p�T�Ge�4�*dtbx���]��+�(��TxJE���~l���� �&�0�PނA���!�Im���>��{���/��A���BLnN��%o��WS���{��I������Ś�w2"�o���=�:��0�eQ��	��"�^�{�~c�=.��/G��eA
%��8���[�eRe�'*�P���+�t�1�f4T�	�W�Ax�T��T0��(ndrM���nv;�Z�L�]H���ck��_�\����� a4|JӔi��3[��"�T�	1�}o�^�'�4)��k�슂xpW���C�*=o������̜�Y�����5���;>��s��b�!�Q���5i� ���Ya�hs��y�}��5��פ�	_S d�f$��]u�<Z��\YJcY�2�A�\�C�ɂ���W7�T�j=��w�H>*�v^�L҆��j4��Z��u�qF��AAI�.x.GŗOrI�`��&�M�;�y��j
 ���
�S�J�i��'�Vf���'E3�X�uŌ�/���������\ju�b7t�8PU�!%������ljQJY�+ֿ��@8�j��L"�o���@�kS���� SZ�a��_��+�x߾�u�ƭ���7��b�ƙ�"�ݬT4)8�@�Nu�J�� ��v��L����Q_��S�0l3�ޮ�9j�p+��4�s-�Zƿq߶f����\3hi�.��	�=6��v��ߌ�QqH%p��aR}�@�v(N%u�>�	P�I�q�����Ji��N3R�3C��\�O�k�1��X��G��(Q�
�e�<��F�[�?�f���Hk��y�

��޲m$Ϸ/����aFJfx�	� O��ӭ%�<��n��mcd>�V�B�X�z�Rj���P7�=�MMF���j6��a#�n�&[�[�Q�]��C�|������^�|�,�
K.�Q�/
�	$*�������G���P��o9?{��?Ȣ��}D<��%�&�X�Q�s4,8�����?O�n̍(Y
��������Akp{��������!Ͳ�_ӷP8��H ��J̽�ɵ�)|���"֊�U�ګ���z�: F����A"�-��S�[DYŬB�G�8�~�8�_�I�~ �MBku
��u�C�	���5C_2H�]��RPXp.�ZR`�ߒP5� ���/\�9{����Q+y�ͶWz]�(#��N�`��'HX!��<�D�7%��@�(�C8������"�=�&�[^�c3�"
-i��gtvP"�u=�iR�.���}�u�Y��0���I����'Q6ە�y��.��������ֱ嵐�$i�U-���g:�RB���A�ΝT=#U:��`��u������p��B\���,A�	�5��L�����*Ihux����O~��8\�ҾĲeJs'hț�t�*�i���^G�����(Ρ{�w�J��%���҄�^�Zr��;���2�ysx�'�Hgm�@�3��NN�3&�Th���-�;��������F�(,{�7ߝ�ÓyX�s`�"��Gd��泖턖�vkb��$���U����\j�<`_#Q�O+x`�Y�RQ���׎�IP�G7��H�<@�9aG�ńH��:�+�<�H�}��� �z����x��Ru�	���'~O��甎��h��(�zը.d�RR���c�O�З٥T���Se�����0��{�ӛn�_�ౘ�M��~�����EeBx�vX��bi'�C1�\n@3�"Q�d�YXv7��w��0=��"�+��Y���c���9u�C1$��"���ך=��]�ol�8�˙fb�(�)Q�V6}Xl�}, %�Y�	b�vz�Z�˧x�W3�c�+@!� G�W�^p@�jp���+X*��!��4�Qe�J���j#������5�53+��В<N��V8����YU�yǎ=��Ā����X+��
׫=;NB�H��<�]6�z|K�q��?��i�NSd���?`q���(,#&]9��ۄ���z�`y�R]���-��#�#�3H	D̲MQ+GM�uo� O��n#r�5Qs	���]-�{0��t�#�.��8�g,ˆ�/����������Fvm����~����R!���O��{_O�[ŜM��T7�(#>E�E(�y�

G�һ�D��L����l�v����Q�j���>b�X�eC��0�q��`�Y? R�H��5����� �<��5���2��^8�0�	�2 �ʹ[. ����J���Y��e�O�ZC~�J��P���NT�`n����0v����0�3��C�V)�m�`;�o��V>���6��пav��������(�8eN3�FG&��,F��S�H�珜-�f�h�r�ן�f���� �C��ȳ��R;�֧Q�IQ�y�RBꥄ��3�a	�f��p�����'���Q�ɲ�o|� �e���N��:]��%sg%���g��OV��n�2�\B	�[�Nv:�� ��I�aן- ���1:
㶠i ԋ��'��c�ɷ���Iҧ������Ӗ�)AЮ4In=�6��6�a�ܨ*��"�5]�&���k7��΄A1�)�NpQ��M�W`����H�9A�8jKaE��/��*�$[��N��.���2�\p:ε	�;�Υ5�.�No���ӧ���I�G����jJ�����s���:�
f۩�;5��xhk��;~�CJ�uJ	�.�p$�J�����<��H�k@>��~Jڱ{��Y��g�r�~��B�hu�VP���0�zʻ��_�q�<lC�{^�pk�:���y�������>C����l��R�����i"^Ny�d��?��5V(�gڵ�G��qw#3;���Lvg��S���NK��1?�-�ؑ�}�_i�n(���h����0M	�lZ>	.EL���w>h�����I��+�'�����;����0��;M�ԢP(��F��G��vx,$��@<�(Zgfu������вY��`�%���6��F �1:��%�z���˕�טq��L(+�˃��D�(��Ej�=�s���ˉ͞N�߈
������عt~'��x����JHu8ș���>b`x�����`���d9VlWq��x��nN�Q�f���$1	E c�am�`�m���\G~�%S����peK[����eJIO�]����������
:�����6}�3G/k�̖�pD���G��gh_��	�x'�����5>�̳O��n?�,7��n1��a���W��!��C��*	����í���(�_e��
5�
Z�L��2���>B!�)�ZC'o1�![i]�����7F�ϣ�c���&����S;�l��
���	,\Bӎ�$��$��||x�����xN�_dO���Z�W�3P��Qv_\��65V����$&�.�J������Oc+s���k�Z��1�QS-6����j���[^����J��EHc }�d�x�N	��"y�_�i�X%m&���T��q\���M��0�	�z���5_ޅ�|�x?���	P�b�[S�����w��"�\��$�jK��\J��j���짣��	�)��ڢ���rS֐�E�|�q��h���oV�+|tp�XM��&+F(cQ��(��HM ���oW�v-��^i8����$#
��R�E�3�댍�������[����K��	��.<&��p�2��/�#!YOw쀘෮�mz���ޱ�����ի�����S��or˴�_�
RY-��]mSa��?AѹYe� �������6�UK.^��ٺ��.��\pD p����Y��g��&�z��k�
O=�#V�������<�s9�%y]��{�́Ĵ{75&��v�Z4�4����7~"��n�O�.�vx��B�0\��.၌0i<���՗>���^>��.���Hlb(/�ʌ���|9�g�Wk�5Hx�PԶ�|!Ő�&��Ԯ%C,l]��ji��qq��4���@F��p�����u��mӍ���=g��d�y)�G���aX���!'�C�?�����z��L� X�9tI^a��T�^��V�@�pJs����neF�r��!6<����X~I[��	A��I���}�jE�r�|��j�/f�'g6�֭;'�R���kü�C|��_����m�c
F��Ϭ�~mo��|ʚ�I�c�D;��Lx� �*�U�z��m��.��Н�"����H��;e��8$�h����4�/y$`��>2s$A?YNY�P���Ů�St��l�H���U��HFT�]ұ\�����A!J�{�r����%�����������WX���KC8�c�!�]�����z}�;�C����,W��il�&H-���$��(�sL�5�bv�����DYh�W̓����`%YV0ؽ�\�dn�
x�=�r(�����*���1dtb��D���L�{����df�q�#�b䦻�ڪ)y�
D���\X>}�>n��D�� ���Ը�h0��_�T!烿ܸj~�c$mF�U̗F^��>�G���Wj��O�V�=�Ū���u
�)HeR9�����B��\�i��J����8�[Ҥ���l-ݓ�՞3���uK�o5)���h�j���aI,�(��&�\5�(z��<Z�:]�A�Z�pmy5w�$clF�����֒��n0Z��"��3]�dd�s0pNr3H�S�1�KJ�`pgB*��B����$�P/���=�5�I��&���g��-�W�$��֭Ju=�0Xܺ�!�"���A��b�X��@$����ؔ�WgR(���j�f>??+$S�韫�9=��S��&�{Ψ z�j����K��SԹ�^�E��ԭ�)Ml�厛V~��H��`��Ɍ��;��N4����	$��;������� _3*��8U:iy���u�?��"SQGyK��Mmȕ��n�I����#�G�1!L�Ke��{�Uh�2�{i.Պ8��B����ۣ�R]�J]L�į�Z����b���_�U�e��G���)�R�<�'���Χ�Xo��8Ky���嵭R�?uk���@v�����{' r��ة*�e9�u��x����2NDÿ���Κ����Xr��= �D�qv�A�L ɞ�)3/�����J��n��n��Z�rT	�>鸘����:U)��o��Ì�����˅D�4���E�v����
d����^@�,�\�>�$�z���6��p�%��s���$�P��&���Ul�hG�Ck�K|9�I2)��0Y!�6g���O�S^ �^��,��/�~�{s=) @��^��ە;��7�`����?�dI:nq}���D�X]�+�|�X�Yb��E��"Y�Atz.�'<��v��������R���)�!S�  �ʼV!O�HK��|k��6y�7��5|h5������H����C�o ��)sMM��Ԋ{Z���g��]g��Ʈ̂?Ԝ!,p"j��Vf�H��B6ʹ�����t�P�&��［�������gdR��o�݄&	D-�69(ap�qY�01/`��?3xȏ���������R�M�� ��%���/x45vOLDa�E��62�ځ�B?�K�L��0�|��W�1졏���}Pz��\g�\�Sz��@�,���0�����\�E"XF���
�2�r�0E���Ӗ�;%�]����uf���ya�|��2wD��g�DJ��ـ�C�߯x������r#a�M���K�~~�H�ԯ���T�6�e�
ŵ�z����q��
�����l�~�������c�Qq�J�Ζ�;P3�h!F�/"���|X]�5E_��g"!B^I�	�8$*ACyS9�̭�D vp3�%���Z)B���Sb���ctH�%)y�8��X��A\9}�ɀ_�'�;\�4�0�֌���ⱊ3�JW�\;���r�"�|�1o���^�lPU�*�,�*C�V� ���"�V������R01�5����e���펚.����繭�O����&.����ш,�\ � ���$Z���k�"��}|r1��g�b�XE*�5�O�#���ꟈS�Y�����7�M�#������r1�=�[F1rF&��0��c��ud�7kag�L�,Ox��r8�����x��4���7O��u~�����`��Xi��iM*��sJo������̔O����2���� E�q��T��(�61+M�c�,φ�]&7;%kfȃt��@��3p�-�]��!4�C\�2�X	���mY��Z��"���pe�ļ��Y2W��'Ƨ.�Yk��ͩk�z�d'CC]���L02�DR�sX�?V٣��%�1����<]�����e��Cu�xo�A��A` ,	��Y�LҀ�_�|-��}Z�Hl0h��&t�8���4=G�lTy:#.������w�� ����GFR�/�;D���'�o8@�a�u����⧺&�X���{N� ��[����2$��a�~��(ʭ{w�������j[��h���un'/��È�a�5��W�\����
��d��ĵvp�,s���h���mB���j]�`����Y�]�(߇��-��*����V���
8n� O6Mh�/>}U���E�8��P�u?ĭ�VC�����y�]ޡ		B��
����I:�����U�[���b�?�a���9�1��@i���]3}^.��%h\�K	i^V����=N���	��%Y 
s8��(����q\�{���Q�H���I����d���)9D�l�,����|i���wF�+#������nGr21���4&�zŹ�v3�5�i@�Ә���k`�#U]�C���@�9���8 ==�!��̨I�H -��8�-4�&�GG}�ܾ19>��pچ�EI�5�8�Z:R�~p�寐?�zsl\\]�|��VTfZ���W��ʑ$�nƨ3+��?��M]K����%qX�٪�Dѓ��w���X�|5T(���3�_��<�E�s�7���ٻ��a�\5����uӝ�C橅ʝ�=�6��#m�t�O|���m����@	"Q��}:�1�M��z��Z�<��ł���*\����e��	�M�Z1QP����I��Q4JGZ	��x�2�I!ƳaQ�GA�{�(�;���! �~��lu�����-~V������
#��a*�^�Fm�����0��1��@�d��9T<xaXR�ۓ��S�K���L�Mi�~o���{b�cqؖ�|;I�)����|;���2������\���yj��r12UQ?@q�������dD��Β�|J�{����/�)�>*T��DܗLD2uA��y�~l1C�c��~�W`�F(�i��>+ �ve�(Č���}�Y���)�K<���f�%�
 ��T�����&v��Gxୃ'E5���N�S�-�)l�;�VE�����q~L�� �De��)������dW(��pz���^ْ���H%�9O��ϛJ�^=�G���e�Y@���?�k�'wÀ�e�'��)t�=5s�������k�ݗK�kۣ��l�',�*l��E}J�p���V(T�j�7�#Di��#���R6p�xwX3/��x�#�c�I��X)I;@��i<�9Z��(,A25lJ����T�"N�➽�gNGV��R���2�no~#&����\��T
���#	��������>�4�6t\�"���f�5��7s�D�ͬb'Ѽb�gs���R���W)�dV�إ�r�����M� �ʢ{{��W�h�=Sl�_��{S�< �w|���:J�����}�^fv�j�'W|����68�C��`��Y�f���c��߿�P���	Nጫ�/��hK�k�12�ZwW�t��ؗ}��d����Ϧ�O��Qf	���V����b-��J���C�*�)N��E?l��)��c�#U@��&���'X��C
�yf�S�H��
w���w'�V��*��������f�H�X8�6�&W���;<�f�s����?���F�o��.o-5Y��i�v�r� �`tRjq���̕#w��Hȣm�M��M�n�:l�L���ƍ�iQ�w~�r�� V !���iXa	���LyK@M�}���mtw}��J�������Hudk=$�Boc@^��#�<�U0{g�C��~AC2/|��F���Ś	�λ��w�S��Ǖ~Y��'O��%�� p�J{�Fc�cJP�;[��C$�D�-�d�z�)m��������+�D��Qhw�]��6r��V��@v$f�T4�eu}d�J0��A�T�4Ǘ�(尀��8��L��ȑKᠽ���)s�z��a�	j�]g�w�\q;X����[æW��R��� 'nQ�4���~|�!��� �&-��dF�竩_w�2˧bE��7=1��a��	
�+��(_q ��@������&z��~��ʤ]f�D1��I�ES�U�i�z�PV�3�]�⇛f�돈
�XM8�I7�-opj�����O� �Kj6p!��L1��NlEV쏈d���b�sc����t�|~=�h�������)��Kz�Es �}Q�{_�:*n|��@�$)��}��Є.������f�ӾY�G���;5�}�������HT���b-����^Uay�z�2�w�<#�}F�������r�C����utHq0�e���7%���厌������=7�U�Z��h��Ɍ���J+���cp��Yĭ�4m�H.������En�>^Q�T�� ���
��@���B!����� �3G�u,̳��v��4��/!��>h �!�"�v
�Q���FY���B@D-f�l�E�w(�V�URR=��:����OG�m¸y���Q:Z��@�pC�>\�=:�����H���sȉ�Bd���;�5[��2�c7"�
�.���jc�M�x�$��p�/�+D�c�J�G&���>�"Y:�A����u#Sգ��1��X���tE{2h�o���;[Qڴ�z�_,�3F�����}u��Dݢ]����DЃ+���U�M	�_��5)~����qSpp��;@��թ�,ܫrI�3�N�zIћk�;� -�i�`��1�D�m��k�3AKûZq�CҬ������m����C���~�#�
(x��"��M�%$��-���}j���P�ƐErRL�Qm0�gz����혿�8���|����H��r�|���oj�*|�]�5d�e<��r�t��ko�Um�Zu��"�-&�I�)�H���49�H��Ƣ��9�SP��Gy,�"ֱ�5}��66���!�g���v�f��[���i���8�@;$	H��>�ct$X�@Z����F���X�o��sZ)ߟ:4!c���x����|iy,�]k3�V��+�q�n!q��os:��vJ��&�Yj�c�?f�͖g����5���~�����*w������>Gi����Ye���Fa�J�YgT�`m'�ܛ��0�g׏H$��5� ��x�3D[���o�0}�4SQ�#>�b�I� �о���}��S�/{S���^���4��V
N�	l5�6J�zWl�����h*��r���G���xH`�l��
�Z�rC�;��6�s��p��V8�Q��1�t��{k���!f���3灒��W��V~����zn���#�g�C���4N ��3��2�͉r��b/��v��Ǧ)S�SP���b ��Lv��r�u��谖%�b ��%���e��{tzו�O1
�2�b�N������D����\B,>��ފ2�j�lYs��H��%lY�KشI|�os��}��+�e����?�s۠w�:J��34�=ۆ�#����kG�6�8��b�੢��a��6c�`�nS��Y�5A�pےO�%��%�$��S��]���iH�v�{Ůr�U�7�g��߻�:��$����Q`Aw�D���l������-~��p!)�.��\���dQz�����|����ˡ��sS1�������G��P���E	b��4��	��:��tL{���]޲�G��o���!�9����uY��᳠b=|~nv��7�qk�W��$-�	�?O��'����	c� @kZ�},+ؔ��l;��	J!����v��V���8��0�o��$��_!j�@��U�����:��c��&����� .#�b<�ฑ�/P գ�X�BI�����m�\~������݉���"��,�u2>BGR^�=����� �B�]i3��g�126�w�&|�U発�`)
������E(��βt��P�+H���ޤ��嘆%�ܮ�>V��U/���qКj��ݨj��=1��D0 Һ��E��a�z����ٵ�<���ߺ����e3��뜕8�����MF�4�fv�$��r^�=p�L��q�(.�C'��0���Ȋp��Pf�z�D?m:��E��:�q�]l����`�{�_F�����䰢I�{����$�բF5��TQ�a��V)�¸��c�=��m8z�|�������Gҳ��{)	'
h}7~)�uI\�se��D^��:����O��(��P�o?��^�1+Ix�ّ'i�*�rS"� U3�p�e��./?9�'a��x@���Rro�rt�C�Ӕ ���)-g�ך��"�����,�HІy�珌;�r��|lޮ&�s*fe���)<�!�b�`�4mAD%k�6�n 2����Ѩ����9�Bo��)���x���3����dN8��/cU��|([:�\""��[���9Btv$%z�^�Z[2��ױ�zð�f�ܸ#�3��r�%��Tl�����KK��~�_=��y�*l!�7N�;
�C�l�kX�;[��_D3[�҉���c�N�ԱuF�`����ߺI1J�C�i9>�A��[��DjZ�9��3��
X)0�E��a�қ�ѵ��ӝz t�7������:Y�Dq�����R�p|�j� ,}����CwmrK04֭k,yC��L�K�#��֖R#(�b��l����}��E��k����f�Q�V!�Q��~�m-J�����:��|�4H~��k�'H��|�_�0���7����O{�W$��z,�Z{�
�+ρ�]� �<�����P:�%�&̖���}>��c�V��Y�4�[�cK�fN��"���hH#͞Ky�1͙��@?��� v��!j�u�$�W%�b�D��o��W��]Vq�5Z�	mx�b�����(�٭�/E��O+�0X��;�P���\Oj@���{�n�i�lp�$+у�]➜J��s�F��g�2x;n�W=*U��)��s�"5?~C�{���;cs(��7I9^��ڥ���߁����`��|�kx�PA�U�"�ʗ���p�[�x��>����e���a���Lz���=�޼�mʀ)�?;huU��z$�Jf� ^�S�k�w:�k�l�����M��+3a�q7�������y����[7�^7�l�"�g�ܧ��G|�h�8�$R��)��h�W8R��%ճ��B�0�F(�F\@�ù�R�����V\�a���%�_9f�F4K'id��qv�g~�/�#�&!��3�]zX�|F��#v}���n�$�� ��COD36q�V�]%۾��_mnh8�	��\E�G�ݩܐ8�T��u�Sٶ+Iu�/���v�k���9��%��2��ĭ���!��~z� @VS���26r��i¡��^��$��ڮw�(��I���B�3	��d���oh�R�p�(�7�ua���=3�2�.�x+i���h�}�Ra����p�c���8�'�#��45��<�G���:8z~L�m_�@�.A���K���W:�,��ӊ[�X�=��0�oe�>������j�G�k�a�����nB/�Z�I��b�'�@�๙�꯱�d�����q�T�~"���g�q�N�]q�<O2���^1��l�Db%��ӳR�����M��myʂ&�t�f�v�G���^��-й�����%4�{qT]GL��g&� �(�6����Zyn��^|��IC������a=�����&|�`��E��uR�<�b�٣~K�P�Vn:��=x����^�l)�$�fF�؇``��ҵ'�˓d���B��1Z��m�"�Ƒ��I�^`�r�!)���>����(	�8<s�i@"������V~�`!v���PU����]���MV��F���ʯ��̔��A!seQ2*�W�J�i��{#��cXq���ư�REh)���GQ��7ڋ����0�)m�������@�03h��Ul�N��χOj�!u_�_(E.`���4�>��2y��'.���ʦn�y���mY�C\k�2�'�� U���l�t�������>-<�@���o%��7=yn���-^��/�q��T(��^Ɣęo��v>:�*���P�ǔEs�[A˳į< � ��SPJ�C��Ȼ�CW�/��hd���o�
c����["�9J�&���'�z�� ���������ԓMJ��5#�� �=�Mȃ��������h:�td@-�;�+&���nx	Vb��� F��jS	^�sZ�$�:_�yR�x\�g�l����*���\�^�3�cGT!��E~��ޥ&=�ڇ{�:�������+	��+�����Ea�4����"rO��TtX`k*ww��1y)���@���4�p4��n���z����=�A�
���u2��lC�:�y����LwK p�ܛ1�ͫ��Y�`���Z�N�=���-�}L�&}���s�N�?ijIB����{~��3�5X��3G�S���D���P����ș��`��X��ЉQS"!��	k��a�9�@+�_��wA#�Sd]z\�x�Ϭċ��L�P���	���M�ȯT��!��x�d=y]��&vЈ���0I�GA���a>��/"��O,���v6����)�t)��P�~i{h�#s�!<-�1�ƙd�A������G҈VQ����@y\A��s}�$/"�v:Bq��G#Rs&-��=�>%�*<N�BfN��d��k�͍�	�{�0E9� �_��Q��M���(,G)��1I�_�#9ê����R��yw�V�{�Xse���Z��R�Ƨ����u)Og��86�Wq~j�P���`ѵ�j��nh.-t�����4!�Ak`�\���NA�~�H��r��$�7��F�WXԽ���jjN�0���2S��t\Sh���6@�Z��dVF��dw�bW���9s��Ll��d�MTS{�������	�;8�c�䮮�j��g�<W�n-뢙!e<��Y���=g�p�0|��{i���ɚq�ֲ��Q L�â�9��|YZ��v�E�Q��y(�~!>1��^Ѣb�[��uQ����Y^���_a`��y�3oT�8��f*�Α�,T��fӣz����۽���~���1��ȯ����'{�Pc�͚�w��!�-ǏP�^�M��h�g������2z��fn��̹�@%x�K�l�WiU�m�$��S��]/u��C�؂���]�
��x������a"ty�&�Q@Z�\\�����z�q 4i	���TIx�����t�%m:5Y��Nn�|^��%�@�`���~c�nrP��[�GF̞e�ca���I����
H�|5m��2�)41K�q�Ee�;̎��I�0�-x�b��:��_�9�o���Ҧ�xj���Sj���Sg�#��m������.[X��tn�8�u]���������w"�20�;+�\��d���E�6[�������kpF����z�����3���Ý�`ϹW�s*��Vi�2H�/=��T��r�yF+��4��4���$"ڨS�f>��q~_��3�9�o��D�L��f�E
�˦5�oˈ���x�wYu��Yk��
�����ސ�ػE�����Q_��V����ծ���;<�K����j�'/����G�H%��K2�w]�YAd*mpO3����]��e)Ma!��cQ;B%₯�׸l�4��|v�*�򸩧�e�-�~�����c��D�j�bsvԴ����QY4q�s�LUD�"�f�|���8��W����'E�~����m$�y��^�.�f����2�:��,s5K� ���R%~��3��w��q��ـ��c`b��'7^���ݲ����ߡ:��)%Z/V���6\�3òC�m��s�'��H��-�M� B_P��u��O'�a�c&�P=�iի�r��^�;��!���M=5i���Mr����(��A�t�%8�������D;���e 3�Ğ����<�u��Xx�# �M�,�7w'����_��4�
�;��ľ�(��}ṃ��4b/�7�g�3gf�E�H;�53��i�r����\��[ImW$������#���8��+ɒ#9w��nT�D��p�p�?q�솷#Ys�/V$L�r���I�MS�m6W?��f�������_���\�iT��>ۢdD�8�'0���9���~ ly�G�����Γ?UX�Z��򮆫 $�g��c��i�$���,3k���K�Pk^l<�}8�K�Y��1 �5W��9y�5��T�H�]�(�È��X��=�q6����\�*a^��o:���k��u=�7/�_>5�g8�ꗻRX�?Bc~�r_��UA�'�7 �)G��������v��eu�9��q��.���Ϸ��͗�ɹ5���� ��HrU�Avu)7QC�U��@NO J�g����兕u J-l�=0����/����ʝ��.�,��N�ώ#D�Ե�|���i�kŏ׮Eo�ɅZ�"eVFNTѥV��M�E^���j����+q>��Jxx�ߟ'�uW+����1�@)ς����a���G����l�����8�c0�O���nA���0��m"�)��:�� �'�Z�+h�� �ҵec�X>���G��K̞���v�"9����.�.,���*�(rn/������?�>�kH����b�bd'2!�B�'�hլ���,/ �'��xg%6�ʙhvc��Γ��{~�($�Y�Ңq\	7�Yj�ô�Q��ѬIN{��s����C�ar��vr�������zDC��K'5'ޥC(®b	gEf�c6�K!B�':�@̺�����t�Y�Ҏ����sļ,aC��>'q�g�8�ʧ���ޠ��+�4pur�1����Y6?	�ï���i א�7�(�[��v��/&:�������ۇ�����W-�����ͻ^��� ���v�ՊW���"=��Q���͡�Y�����2�d���|��,�qH��#�C�1�o܀LG�����2���ۻz�RZT����A�bգJ���aB�[���V�L��X�S����x��.�vڲ��65n=Z�޺����HIN��ǽ�~;�H�]����;�<h�@K)8Y2^�1�������i���xQ�Bk0�ME1�i��Y��,{5�ޮ�ss߉��0Η�z�&6���Z(��K /V�Đ�f�eJ3*�r*�� +�L��{Y�=F�Y%�P�*�Tbt�n���./5���t^���r�];�Z[�
^p}t��]�D�)�h?�Z���(V.܇������Ǳ�������#}h�X���yk�*�֐dX4�<J�0l�/���'�����^�1OS���=bc�c��Lar�v-c����X5FO�5�'���w��YO�w�M��{�ŕ|I@�ݱbO�J,��I�����8���M����Y@���#�܏=�	�����S=�5؃��N� �S��ٗ}= ҧ�p�ã,��BϢ�ni$.�t�Egp�B�Ie�d�������Fr�	u,Cm�B`��'"P��uK�kq�9Ѭ������e��Db�	Bm�'&��*.�R���kP�o�g�"f��4KYm22PWdv3�n�|��z��s�,r��@h��ےP�А�a���Prg��n@�
/���������Q�L��+�~tB�m��/>��%�����F��~5˦��j�����Ϥ���+��=E��2r���;�J��4ܨ��i ����!��gK\8��q����^0�g]��m��}~�oa��^R��R�,��$��R�F�0������Y1F8�س�N5+�B�B 
��b�k�:�#����Fd��g}�^��UD)sfS�����^����1I�V�v�c~����~��Mq�&���#f~Q�d�"���%�L�J�Jڊ1�XX����m��feQ]�jҘ��R'�}�g�I�b��\�(a^�Lëb�8�65/|��78���T�pJ/��z��3����˳��6��<RL0���fz|1@J�w�FR��7��]�*!�6�Ϯ�q2�7�(q5g>&�o�U.�����U��&���##��.4�Ki�B������E�)���g��!z-�7�@X�SHm{�v����������L{	�6P~�57qn��`s�������6_��{���[���F-�M�K��Fm@���Cl��[�d�%Wa����NL�"�B�ɦ_�rQD�ɿ+%��ȷ���ÒWlM�t��@4�-^7vVX�7M��NS��w�ڀ�q���0Dr�l��3��.�H�ݷ�,��g������z5C��h3d�=^9V� n="0h �k�^1���M*3"Wؑ�Ħ�"�NE��c\�B�V-Wgv������lkg�n�Q��Sc/�pٍ+4|��u�fR@��[k'NAl�� I}�b( 5���
6=��2dǻ�
n��sǼ���"����0�hsCITj���͑^6ƴ�ߟ@ Ǣ���W?�)��?�%/�9m`j�4��}}��k�.�V<��d�j�mӪ{��PE_E����ᐈ�>)�я��_�Y��q�q5C��_P��RO�!R�� 󾦓V���rJ~O�u���Y�j���k�s�nPf����(~��ƼC 0�D}j�Y�5*7��Ð�[�hС�䚖����ԍs3>g".���#Fo�ŠX���ltǻ����'�ݢ�;Z�g���y*�\�=)U�JyU�w������Kh!����U���N����.���:�7Ĕ���.�뵘p�#����~�D�^���e��vv��\3�W�/��_sC�ɞ�?�j��:D���r���&�Mt+D�Sc>�e�� ���Z�Cʊ���I�d�C��z�h!�a�@/ݞ�0�d�FT���� �q��#.7�e��TC�F�wK؃����o�0��Q��g���y�b���K~r`���4�5�9=��t�����Mr��G񣂓��	�oO��k�����\!r�}y��u���'4�fI��^��.�.E�/�4'wڸ4�i�.�`E�Ή����EW�\��*t�XMò�Pc�p^l~cYy�=/�XL��:�r-Gt�r;��lʆV�B ��VE������*]i�}���o�O�V,)jM���d�OV�H��a���&87����U��>௬��Ǝ�0��ۺt 5]n{�]7��0h�Sl�9�o�F���w����R�,v��^۝��T%c-���&�;���J�V�ω������K�F�Gw����N�>��^?xF�b�F�ARu(�`�\D .�~RjVL��q��ڸ^��{o���²ۡ]ސѢ��{�X-�9�6k˹�6+�ţ�J�8�n��B�I�WE�(������dq��k"�����d�q�ǽ[��MS�������&[~b4�Z"8��6�V��!�2��R�&��D��d[R��������l�����!/�k�Oс��9(en�%��:u��T ��I�i8;~2���������JY?Y�l�����x���]���be|�̋E�"u��e��[�}���ןI�P�q����QЅ\M)8'^T�,�R�� �:�ˎF��qH��1�|��9[,�M��'8m5!�g\XX��	�$�E��t\�#=��+Cac�&�Ǣ�YYNg�q,�Mo	(?B����	ؕ)b4�g�¶����V =0R�B�;0�->,��PxM�O�
�
�Õ���vMɍ�7g�6���[E*2+���u,8�8��`12�r�Q�ь��bfܫsN�d�B��n"�.�+p��8����+�}E�M���U�$Dt��>g@S\��q��E1���]B���`���S`��0��,h���,\�(p?�M|7�F���^�S��Ne����+M�½7����_�=���].=�Mx�x*��M�K�W��6�y
���%����v˒���U}�ads2��`�	�}�L��!�ţD`KIe�׉�m�S#���Eт+��rYjf�T�xkR
+&C�~P�Xi�7��� p{��j��ۤ�'�
jo�c��Ņ�$�xG�0̔�I8��h(��0M%�)��Rh��]k�r�a�Z����s�CqiPT^7�5���ꪙ��oR'}r��j�o��L9ґ]�",�˾P���K����%��a^:.#Ԇ�)N�r�E�������ҧ��v�5O9`ɏ���֚��H�b�u�*��X��[派V:\{6�N���(*��v�:=*�����78U>� ��7�7��9	-`�˻��*�A����ȼZ/X��e�4�a�2%��T_����m���B�ņ,JR<�a��Fp�D���~��'zm.�64�(�Dn\(^ؚk���5��Ġ���zA�H�9��F�#<�'RA��^XG�j��� y�7���ڈ�.� sa�t���_MT��ڐ��s���b�i�r�_�?3�L $,i ]LT=�"5s[����?G@��)|������6�O։�Y�� ��a���]���8q�'O��2i"n�l3D���^�&��<vy0�y$J�\��%s_e���»�L-Gt��}^V���i�d �;�*���~�h�9#H�f���`���'^�Z�B�3y�v)a�F�0QM�&nPԌ�J:�36�H�%"��U�؈Z���40�kgY��4�#p��u�*��%�LZ7 ����B���#=R@q%������G'��kj�S��l]��	@�ä��C�"ػ�{0�8���6P/�0Ѵ����ʕ&���:�c��ܫ�zI\�B;���� 7��1B�FԤ��M�R�x��_	��Idp:v�
=W���|x*\3O��\H=�l��_�Ń3�5=���2�ɯ�PU4Ls�������"s~;�:�P�@!T��=S���TH}�r�2A��[�`�(�����x�"�yބ�����A���g��}��~-�N�p<�-�J�Ajg�.3�P��D��������q��1,~��
E���</��Ԥ� v�^��:�8V��mp˽��>�{R�9��9Q�c�L_��䤡����6(�6�'�*�'#Y�P?���"&���7�:���@|��Н�	����j���ڸB����B;
�T�Ȕ�/�w��	�]� ��F�Q��LJ�¯\��|!ω��v�c��4���A�����5��]�S�����w�QڥZ`4 ��B�Y�"B�~��
<uQ��#&~���Z��2�޽t)�@\jt�r ��_/�ږc�O��� �z5J��� ^+ӻ�u�]���~k��E;;�?�\�[7��=]hق��IK�����]�M����MwY��yU�YK	� a _?�v6zvwWK���E����c�R���ݾB��vH�)Hi���!�Z�Yg�׫�H�"0P,��� RV��tp>�M~�g8�˨��n���r�ƙ�XV!q@��u�;���e���^���;�r����Q�؉��uL��PUl��oVȢmcCVZ�MpԷɹ��C�'-�3�٢e�E�t�K��%��sՕ�a�� �00���:���X`�-�f�:F����V|7��EZ��	�P�C���U=ԝ]�_����6a�f?F���h�YǶ^s�r�;�2�����Vz22�q��R�N�Ss`1�36dC�-�؅���4��Z�<(if��vD�n��3�7�M���w��u��n(E|L/���t��;�VMJG��
�k���!��������-=:�vǫ�&֣gxM�����C�2*�:���Z4�2���M�a;y��F�ޛ�H;��Ԗ3�p��ɕ��;^c�����3�WbM�I��(����9V�\�j�*���;nmëK7�m�-�M�z����K��T���=$���꫱N�c��od�5?�O�m-(�Q __1��f����B��ˎ�:�겨Kg~j]d�S��M_��3���=;�x{)����Q���Y���*0��X�_W�/� �}Wx�:��J`�"���+�#l���\�;1:{��վ��;�	�)���2��tC� x����!�R�~((�S��Ie`3��5�	�,'��Jk
��0MZ|�9���C]�,���`�a#�����-!k�N�R��D�Dh�$��ub*�����Qϥ�
��3Cp�n�?�%T�ͺx[hy�'7�ٍ´��6��� �ۏ�gq�H�/��M�"E�<���u��y)Rf�4d-�΃�f-��8k�E�9���*R�Gz��~�x�Ў��P�%����/�g"w(��nF�;{Eӡ�T��6#U�Ž�/���CnT]Py/{n�X_�Fnc�ɣ�'i� |��rp|�V0\l���f�a�������;��,�y�|��*��x�c�
� ��^�ߤ�gAR�v:�r���[�����<>�&䗨#�QiGдi
k�[��~�Ӫ5r��M
�6���^�-	FdVOKHQ��tiL'~������^��7KTn8J;}�U7���'��Ӂ�Q�U���������L�~��tS�.N[��c�����"��}�������w"��`�M���l�+����;@��o�!��7w���R�0���*�<�-��9���RgI�.�%�-��z�5��J����(���"��,�i�i �;�欐�\JaJ_**Yy�� C�$����p
����. m�)?�f��� )c��F?%7��C�����W, %+dc�	�1wS��a*r}澆�k�����:���.�)h����z%���J�70��P�($HG���������E�_i��48]v�~��b���q�,>�S�`
Z#4/� ��۵	�Zḣ���e{��P$���Z��&�Xg�b��݌��p��Gyh�� ��wnO�ˈ�>e�s)��a��T;�y��#��^[t�F��45����K�����`/�Z���S3�7���	GH��ٻ:���x�Uәꁨ�i�_0>�	��S� &R����̥U���]�H����,
�կ^/O}S��w����L�P�����[��݀d�LV0�	��q����I��J���m�N�ģ���g�^ڎ˔�88T,���DiN dP�߇"/�$�׫�Ʉ�rm��׮t/p��-��Nu�-5�6(�v ������jLvVhLgLV�yK�!j�¬~�u���9S�*K77��Q�=gq!�Q�f����+&s�G�:�K��B��s�'�"큯Ȗ�̊�;ƧF8}�Ev彂 �p����[�}|jȮU4`�,6�r�M������'�|ԚPx-�_�t�(����9%`3��K{s�q�b=:�P�k�}ц<J�
/��W�n	�'6 ���A� H���f�/�C�Ԙ+��d? DN?�����޻'��%V�^N�Љ�(:�1w��i8�R��B���@�&������d����'��S/�-,y��)�*������y>�
7�>���K;��H �����N�ݎ�2_>r޴x�|m��׺:�I�/��Ȃ�5��H�pN�j�iP���OO�(��#����WAy�z9�����t<@����"�Ԫy��M��O�.m�qO E�C(q�Y�;���C'h�Rc���'�R��a�s59֠�X9���Q�Vr�^�$N��dט�9���21�[���t��3�w�$tolR�����c\Qҝ�x͍�����18Δk@>�"{�A#
<*�D�P��@���+�� 
�\�
5u3x?�"kb�clj�'�M�	 �6��l�0a2��jd�L3q쮄!�x8��P56���FQԭ	"�0�N�\
�&,d�uox|�̈�}�+N;�ɗ��o!G�8�h0�#Q"��zɉ�s��&9���O1x?���k�\V-��B���n�����2N�r!�B�.He&W�M�H���M�)(|oF�x}��'��Z��>���dk� p8�{+�9��/�b�PY6��r��$�Ie�#4�.�9��N�8����^�F�M�@�"����*�Ez�Е �&�iV�"ªk��q�dTp����*5{��N�ԧ�}٘���WW`S�%�я�����4�LI����j*����;����0���t�ycƋ�=M�����ϲBm^*4�gw�T,ڨ�8�K���l��[�&<Oe%�Z'���(Å�)�Wv��q+��n��-���!�'K�\H7������<?�����e����G��(6uIEM�C��gL�i�t�`���u��+��r)*�'0���#�!|}G ?��?��ۍ�:��"~%��
�uG]�־���V%{ڀI*[1�R4�PWLܧ��iU���������,
���$�3}?������к������p�������a@I��-iR���_� \02\����c�־����"]�œ3>% /Hj��Y��4@%��)a�,����%C�5#�U�b�f��,�j9���̈́���rm�@���U����cK��/py�)�n��'�a�p����l!�#��aHw�VBo�����~ɹ/��K'���Cիe:�Ӿ�%4#�����0�D�=,[��� ��OҘZ/�Y�]i��+)ON��(�멘|N�C��f�Ċn`�▩^��u�~�Fu���yY�XbOg�Z؃�W��u����gi0R�x�_�J3Va��.)ON�f�zT�N�K'��SH��bh�1>�tT+�ČA6��|������ziGe�q��<4�-5���[����@�
�S��_���x����HY��?������� ���q�D�	@)e��s	������3H)ğ�ܷ��nXy�u�퓭c.�;�iOw��c⤿����n-�vyA�Q��R ?���G,��iG���A��#C�'(Ux v���52~�j��f��Dp�L�� �S �&hp�Ҝ���n�s���J�,���⚒�1���}a�m!��
���7�o��D�C��$En��^Q��HT
-�{��<�F�Q����:_���fl��&Q@#��DJ�1 �~P�}�T�p�}���\�{e~3|>g>�(�=��e$\��T�e���/����*���C�vu��3F���\�&?�K�;���-pX�6���h�F�k��Z��p).z�m����ę|�y)(�XmZ�pL=z�a��.!lb�d^B�L5�#�9�Y&[�%�L�yXd4v:�;������wҟ�Y�"�ؼ�R
vs��w�����6K9{!�����7a��{G*�<�c� OJ��NIdx0:'�+n�#K_#ȟ7��,��=V�{*A[~ic��b���.�Q��>��p*�M�3��0]D�l��g3W�+�e�Om�NKO��d 2��G�R�ݝ�VUN�	&\L"Ϳ�D�H1��!�@�u��#&�Ah��Q�uڨ2�w��ģYڰ?���㮈����g��;�;
B����"�l9�=u行}�^��kBB����G'�����lvo>��ק�E��_��+�X |M� �㒮�,kK��7�ϝ�C8,��&>��w��T�04T������c� ���W��ru�|��$dG�Z����PxP��.E�6��SEƊ���:�Q5E�'�K�'��a�y��`��LCZB��Q��}� ��:��������|7SU_uK���n�!5r=A�c�^�/��f���4�h�=��>�J#�����3�����=��_�Sདྷ-!�[H�BC�0�Pf�HNQ�DH6�DF>���qM����sBIXGv�.gA������e?)���K@�z�lp��섩��W\�b��/��jIi C$&Sֈ�jNc�HeD��f:����י#qY���7�a�X���ie�W�+`R2������t	~p���9�]~!���"Ab����VS�t��`Q{qO۱D�	'��FlE6%_nv1��E�r����z�x�����x4}��8-��Ʀ_�7'�l���H͇�?����17ذ�yo�t�3p�|��gV��SQkͣ�WCJ=/�o[�4��{�����:0�V?����QsM��Ϧiy���2L��iU�Ա�WaH�C��m�X7�����K�$�X�}��L�Y���-%�82e"�d�c?�)�&����͇��E��齴�j᠉����?}o6�n�z����Rep�j�\0�������Fo��7S�m�Į^�C?)W��M���x�ڣH��Q '��_�RSx�%�T?��B�{�\��JlI�u��tJ*q-q�KQ�;�5�!�2�Fz|�̅Ȱϩ�ݧ���*o�n�1������T�U�hm�<䙺�$պjU5���0m���:�V�q�����SO���3+��k��t?��,g۔���S�p�n����;r�a˾<\��䡵uVJ��1���i7��/�^"���J��?����FqB�g��F�B�'+@�iJ�fE����L܄�u(5���eIR���)��m����&ue5~�f�sV(�ؐ�1�?���	iL�b�f"	�p1�#u|9 ������&A#��=4hqM��yR�!t���uުI�9�u�:P�o�Mna�8�9 C����U�?���BLǸq����ic/�dt�*�O?���k�
.��vڦ7mǕ_�L�R���[�
�v�۳Z�-�5[���������/���q�xx��?����a�j�b����*�0�iC�0��i|�c����l���| �k�D �n�Ph6�<���d��m���Ƕk`3��%ׯU��|�L��u{B���y�C��U�j��>?CsK��Y�Q5�>J���7'CN��9�,_�.�[M1�NV"�[2�K�$#W/*�J-�z��\�e�`�)��vg�h�=��+�9����j�2AV v<	b�k:��	��� x�jUv�xM=ϋx�wճcl�t#�]�(��^6cR���S�s	�:ɦ��tW���,>�Y�p�]�M���] �зzb���>��=�+��a>�o�P�(�L�Ǵ��4�)H,ܡ���$/b/,wl_5M!]O_oE�%y?��h�A���\}���P�B�̅Iܫr!��<�tdz���cԳN����lu�����S%p�
�����|���Us�*ܒL�����F:�e��A��\ٮLS��{k� ?�$Z����3�~��
imr"�"�ͧ�wC������n��=T��bs���A^����rQ�E*+�jC8�c��:��F��A��]�}�;t8�ŨJ!��/hu��g�r��T{���Y�k���\�P�<����ӭ}f<0/��V� /J��c�G�'�c�@� �	��o)>d�?p�X����3C��T����<3���+x���\��ţ�{�� ����E	j�H���{Da��qptw ���G/>� iC���	L�N����+a�Ƨ���8t����^#]3�	|�^D����'�x���ʳ�j�.x0ØDw�>�n(q�����ۇNl(� mL�os�g���gî'�5�1nh
b�N�'w���F魮Ѧ9S�W�}�M;.*)��q���ƛ���e����.��4�͟a��5M���`M���F8��Zۣzeq����R��'� '1�������F�O@4�$z]}켝��18n��rg$�#��v;���Qw��O	�̇�fF����b���d.��<~İ��mxԱ��d�N�#hI����p��<��C�J?��3 oX$��]@m�nK��78��@�mqT�����8,M\y;�!MaJ���zt���'o���*1k�'~���Z���'��h��/�_R�*�:�@V6�{ui���i��-�����y�H���	�֔�>���NQ�R!<(d<�+�L�M���rQ4+	��sބ_Z�N��:7T��*a�&J{K�E�Fnf��~��Y���c�c�m�~�A�R����,�F�D��Fp���G*6P�C`�^�dR!@��!'iC���SVk���H;.F���}����=>�BY��ØBr�� ��QM5����цN3���5!�=�j�[�ûxi�.�� U���I@T�|������8���Pd�l�2u3��{��r�+�]��K��fX�%�xT�IL��|�Oʎ��p�M�Ei�8�E��/���J�x����^�B�]_�t�a"�*�p��q��ң�5�t:.��� ���!%zM@t�A�i���S���e��5�h�$�WG�b�N����)(g`v�}�9N����'x���Nm:.�����wv�* �º�S��Q��d^�G�@���%'���)I�,��zy��cǖ�1���dT�Oj������L"
�ᛷُRn�(f(�&���:�l�\�)����^���Y%�UP�ja�Z��M�{}y(0���%�Y);Ed`��_���Yú?����P���~W:9��;O�m�InOVL�7��@��b�K��$��]&�mu��C��"'~��k���P���=�5�FyL��{#�ť�E��ͳ7���0���?DGV����2U�;Ht�o�Yu�+y�9H?��g���c։T)��=a{*�ST��2L�6���w�aj�4�|�m��� ����	7۽O�}Ea�x�c�h�>�~@�$��dʒ%a���A5�8|@]�T��!wW�@�/F3Oř���u��C��������l�4����bEwPw�Ibo��IlR��Ν?2�ǐ����{Mv�ѡD���!���O�/f/�<�{/w��ˡ=+Tk���S��Q� ���kiñlb���4G/R	��f��`���e���	�y���CV�a�m�~gPXou��gG�p}ߝ#U���T؁��l�FQQ)_��_	8��g���ϙ��a}I����#)�"')���GG�����$ף/e���5u�>�GO�e6NT��!A1'M&����l�[!]D�6��,��7�őaL
n���8���$��9�Vi�(yG ���+�n��-�Y�KM��5߾����H7�_����R�+\lCN���0�)��6�-qT��#��@���BbE��c'9�=����n��$R���� ź��2�%�OWrp)� ��W*�?�9��]0��{L�z�-���D%�A|�-#�mxHi��+�m�����^�?�����+��G���4k{h�Aݮ@F��U�]i��0�U6�f�xŀ���� �,ն�A� ����~�A.�J�MWv�h71��w����#��~���[����o+/�Y��qMﴜt&|a-����d�Z�^���ظN��hF�S��V&�2�~��ܡ	ʆ�˨}%����ܰ�����{�����$�	��<'�Z�u��G'h��<܏��(�h��?��h�}JM)
��$�а���T "�oG���Pb��P1o���Ij��!?�&�O�$�}����:�5.)�C�[��M�|�VG	�r���&I>���(�ͱ Ȯ��.y��hb��Cٚ�)��F��������x�~㩿����}�y��l�.��wl�����W�,xYZBx�Mv�T�L�}�?K1�����,
���I��<7I�]��T:���a��
�C�Y��;/<��)V뵩�b&���nW���ri.��� ��DWD�����MJ�4���E���!õJ�CuwGwb��
_����6� T��J�����9H��.�f�f��~:��!"���ʮ{,/�Z���,7�[�z��ľI���|�o�7��C1���V��H/&썖�H�3x&��l��1�e�CVujW�,O�m�ִ��"��	�Iȷo#$�.��¦yF�8���[\�%����y�S~F<m��f
c�dH�bEb�zqDG*�@����eɛ�_Bz�̀{7V��.��*�a;Ē��D��PM�_��4�89�!�K20��&-�jY��*��^ï �/n≓��ݤ�\e�V����m9�h��e�a�|��X�K�H \Þ�tPC���?�c�n�_<�W5׃XF���H����\ I�E� �[��(�6$'�p�RNn��݃��a��7�}o��$�?�a�fn�%M�%J�y�r��
�PMڹ?�p|��p��wu�twP�,L��_�7�MMx��X��#�J��0� ��Cn{�!����n�[h��L�ޞ��Y'.����^�.�c�.��U���7~,&�\Z�h������A�0������P�����n/��4P��ڻ���X�g���������bH|um�샾\�\8�Q*�w�is��Œ�o��Y�NF�5��Q']>xߪl�s�
h-^u��Ɣ�����m�g�2�v�y�dߤ�Ζ؄>+A�&Ǉ��ł��鿻A�ݡ�|�*]�z��4��m�򹗯=P�epx�S�o�����Wm���I��r4��;�Ŝ�O߬�]���Q?cc�d�����f��� ~�[�f$��p�j��|T�7����1�-�_߮y�){B�����
�|>�9K�Ie�Sӷ k���`��U}�$�A��L0�	�&�䕌:�a��g�
��N�k�#���q��z��#�O��<_"<r��5pLX\���|K&�1�RDg�*��E�ȒG���:�a%yj�g�����e�[�*3a�b��n��(�;x{^8.w*��SG�R*����u)x�#�3������ʜ�v�-U��*1�����oec�nx�B�����䑡ޯ�1w\(R��L����g�,���5��@,%s���a��p#�u�D�S��Im��HHo!���ZCE�L�-�LnC;H�|��%?_2��w+㋊��G���Մ���$��ss��m��' �ʓ 9Po��q�)�r�u>ܖ����e�Q�-P�� ����(�Uo<�Lh�s�)��A�d4;z�,��56*M߄b�@�N��{�?�溺W�\J0D���om�xd�YO�����q^���C�#0v�L�!�:��
�=���-�1��X4,[��`���A8�멧�FNf�<V86�{���;$�~N��d����2����6\�� *��ԗq�E����BWt�vR�G-�_>�{���^p	n�K(aS�:�@�Nr��W댯!��@O��Jm�Q���$���'�`���*�>bi Q&��+,O
"��Bn��1dq�SЉBOz������˕4�vV���T��ݓ���'��i¨�@h�t=��@�e�Bi�������"~V!�umy�tքpҕ����:���<��y]�� �w���f)����CN�)���W2驕�����aL���H��L
v7�B*�Ư>���9�z�&�4ЂI]�ig�=�0Z!�tb�S�,�ʀ"�]�Ք������z�lƾm�ڀY��{���[�����$f��Q䉲���`�6tÛ��4���C{7����ʹ��z0(���mI}�g�>�R�\�#�̦@��P~�8 �M��	�\$�ڍ#y�&�u�����	݋�M�_0&?M�_����V=Q*(����x�0�8�zB�tH��$����̜�h�S�b�5�Ru�X�m�]�4�τv��g?�hH���|Gr�ɠ]!�R\{�z��,��+#�r�?��0tN&I���t�2�1����/����B�=`|����&P�%8�??A��9;��}G9�b�u�Vx����?nJ�	��j��y�np�j�#�l�K����<�l��[8H���ʏ*4"�@j��vP� L�qBt��9B��<�3H����Ϧ�Z�q!�/4�P���쁬�c۬{=�^��}? �L��ٲm�z������u��*�ꓵ��>(��e��A�K->���mxT���`��h�Sd��a$A�>&�'����!'�s��n��l�J�+i섽-������ڎ��R  ��⍲J�y��ui>�^M�p�;�d�҇�ͿF���ll�7o�8R���I��؀��X��m��3+m�0=��z�N �?V�mu&�8���N@½�RT���y� ��I��b%or�	�3D�ӓ��j�!��ԟL�M���w~*xY�]{ $4�o������H�ȟ���=f I��O��?�J� �oJTxҽ�r\�
�2�l!��c�V�p`�.8AB!��p��J:n��� �'*�F��T�̕x4Bq�9e��4���ꁠ�:�B��� M�s�ҳ�+�d�Y���9ê'�݀��kS��9���G���r- �����8�{F:& h�/Γ+ɗ���`�#{��I\���@U��F��xԑ��"L�2�&��f�)a�G 3���������}o�=g�vF���rei޿����N���Kѣ�TB����2��M�O�ɗOP�`�	��.X�rQ��.U��i�''e "K~���2���u<A?}�R6J���ɢ 2�ӣ���Q�lP<)1�/�����/z^ ���M<�ȉ�b0�K��v�U�@�nQ��{���yN-�84�5��po{�I�4�/8����1�PVL�谇�~!���׫�Ou���PS�
��V���������~�F�}��ۇ�ey�:Q7S���Ds�����=3_��}�� Xä�N޸��+bK���IfD���:r�ՙ �%�M��,+�5���g2�cA��s�o��U�nӺ�nnp�4O�|J(�����۸g��}#��b�����b�	n����j�ɜ�s5�-|(~���b^�@��hz�A;oյ�����Ӹ&���	|�.l�A](����U�_�pÂ�~��͑�֛��;�,M�"i����k'(D�3�����%'�AyBfv��b����4�J{�4@�V,q��aI��ՠ��8��7�Q��U�r��}YK���~pO��t�����5����V�mL������/��lH�L4f��>g%�M��˼E��펦�4V���*4�a1� �.M�<JUr���͙ ���EːB2���-��ߝ�g�uo�!�t����ґ �t<�q6Fmڦ���E77������J�Nb��f�ؖ��B�)��Vb�mzK�A��]Ǭ��b��s�P�I��.bG�|i�ޡ��� T����wt	*M����(�*�E���[Z߃��?9��3�%?�+h���0��)�J�bݶ9+B���&q����a�
7���u����U<Sw�H�%�1�\'���UN1�����!�0e+'��l��c�EYć�����i6��qm=��yO��f0�I�Uoa�n6i	��ɫ�L�܁��wժ����]�%��:����q��!�c -4��S �&l�Y1��P?^f3m�ۡ4P}\�m�M����u8j_]9�«�/=�:�"����$�j-���>[�����4}��v�5$�a_�MX���[�#��!|0��А��HO���_�]�/D�^��*���6 CF�U�+��tF�p�Of4�M?����<o�	"e�m�d���ؘ����e2��q���"=��ۚr�<���Bp5������Ywq�=�1�.,��n�A���Q� c�~}���9�E�����%�{�\�G�j�'�bN�A#~p�c><w�m��2;��΅����v�q����	��/ho�Qjd�1���dM3�X�5+sZ���"^D�G�YR��|yț�����%�|�a�+^��^YF�rz�ZFX�7�8$��q�n(�X����A��}u�v����9��qRF��qj��4�I�(5Ɩ�I��� ʤu�u�W�����
ɀ=JI������[u��T�K 
���y
�z�,�L��z�	z��SY��9�	E�A��Ml�[�� �(`�l4kZ��;@Oq
c�	.���P	��`\�x���do���`{�
��0�����[���Աq��� �s��D��2՗Ϩ
��DoÃ�$� ȾyyZX�\^��~\�,���j�ɺq~�`����k�Z��mD0"�@'���H���=�Y�l	孎���)����B�y<��G�X�CW�6�Z����q'
�+�ٗY.�F�2����2�ȉ<��B1�x�ONRw�������ƭ�KJ2j�
`�{"�cͰ"���J��VR���z��Q6�q��	�� I�`]������3�ٳ-p�<}]�W��2�A��el�-�y뫁+���H����g����`����pS�9������B9%�вg����ZE���bM��y�:n����@0h���\�����"�w�|���\g��7	䳳�WF���D�,ToڗD�@�ge|�"�8-��\���6>�`���֨��|Q�ܑWXV-~ĳ�t 8��kp�&�i^�a�iFI��1��܂���\��O����Wj�4���l��*%�{����?����o3��-r��5����38œD�v�c~ъ؋6����B)�"�{,�Jx�Ǯ=����g�⪿&��(�l*T�����jQ���;_8 �J�<^��4p���ʟꢞ�����Bko�=B��~}�\d�3R����S��u"�D#l[�[ �OGs27+�y��σ���z��i�l��%@Aċ@(M�v_Mp�v��Oڇ1Bpz�}�9��a���M	�FRYHs���T �m��vu��b�f���>�]��:���ͯΡ�4��j�$�f脪$e�ݼ�:~|~�9��"�rx\�=:��l���A����Z�ٛ@��P�ٝ�'�5�6�|�Q*2I�_��,:O����(8�)��4�/��Mg�b�5�K0�݁xeU=�����wI�?�y�q(��S�C�P���_��b˂I�d7��6|J(�������w/�������c0���$����V�;��LL =�d{G�������Z���E������8��5���I�N�l-֯��z��_d�I&u0E��s���^V��Ŕ�^��$)��?=�c�U���͙y��r3�g0���/M���Z��+��U���(��:�����ԛgϢ� �4����ӟ5����fW�S��8(�T�
�ę�w����%7���M<�	I�ek�k�j#}X��^����K�4s*5��P��"P%-��wy���%���܌��w�>����ߙsu�$2�3����1�`�K����?]ɷҘ���lx�e�#���{�/����x��?Ҋ%�(�"*�ʪ2}�d0���\Z�Lɯ��g��̷�SZ��`��;����R�>w�z�7�8���� &Ҩ�ɴ���� y���qE�qz�K^~��W#��/����'�7/L���<����â%Ib�$���%��93�lމ�\F����D�r� X��� ���C	��p֤���,;4��Ȗ;aI:�\ʰ4	U�s��6�Z���0}���f�p�@��j��(APjB�� ���R��<鄩�#��]�k��(�B48��d�$=�s��4�1D��yP��|Z�4�8�7+���~�8���/��q>-�b��K)��U($>Bi�&ۓ>�,����H�B��a�� 랓�Q�v�-$v	���~|�Y0��o��B��iɛ�4Ӽ��ѹw�+�`=�&/�h��5������&�#��W�R� VH�`1m�4
-�}~�À��W[��`��q�?��9�*�[>C��2�wS�e�#���?(Hy_v���5��j�A��&����B=7�E�_�gB*�K�&�ƴ�6�+����lwG1S�/pk�?s�Wnb,l[������I5���{�g�ݾ�K�nmx#�@�!-Yy�g����o݄WO��3�07���G ��oI%v��gF�S�ET �øG���^A��9(AI�8��?�$�b��#�Ȧ��~�4�drR�k��-v"T\�5PLY�U��Kt%CM����풩,���!�bo��nI�T@�q#
MG� G�����_K����o(��|��B �JYlcWգ~ $�
ym�Qh'Ǘrfd_+m?+�թͪ�hP$)�Z �����i�N�ƼLՂ]�&�_0�j�j��6��&�NB���+L�m��g��a+�n��CHEg���I��io?�Ůf��H� ݡ��!�Z�m������{�RC�Z��L�����PQS��m{A+��������� D̘T��U3�bi ģC�J[���-��~E�$q�+	��Ь\�W51|:�f1C'm�	�"��\���CA$�&���8"pi�R���
���U�.�Ej�~�����di�v^�@y�ke cK�@���%���j���� �s�86 9��|�1�8+�{����MC�=ce�~m���z�4��%<!����:"R߇'��|����?y�ƍ����H��5po��*P����V�<�Ia�S��7����>C��jً��rf�N��a񕗧s��+�f"���Bg������Zn�ׂ���>����%���"dV�|�x���v(�� t�w?�<��G���oS���тs�t�vD�^T�K8=4]�}`T�gW�������q��E����E㞡�:V�����(pe(�퍴H����}�ՊkS�僳 ��)�k��_�7+���'r�����T�*H��!��yV�8���A��&���6���H���\�#��'��fa�����~BE;*:��8��oO�f�i���ѓ�M�(��^�ã���׿}���}���E4"�9;�BTToV�h,�� �	�Z���b��PM�h)B�_��[{_E��h���w�$��W�Wp&of� rtI���F���f�S�@�ȣD�G:\;�.LU��6�R(^�PBLg�Fh:
�P{�5�0ڿD.<�V���!��xj
8����}�7Ř��a�:�;�L�f�d�X�"��##�S5�K*N�}�N�]�T���t��O�_r+/[~PA���s"H��l�g�.���o��٥%���ɴpԼ��3}0eR��MS,1,�3<y�a5'�)gBxt���g���7%;h��6 : �'�Y�L0�p��|��*M +��b��:�\TF���7�ޤ��$+Xk��2>�pP� l/Nn�*]�s��ē?��s�dp�3F�2c��W��vU8s�U��O.�T��@G4��6D%c{�U{ w�*{ܣ=�9�������D�ȁ �Ң:�*ۧb����K�s(��b��	�f)�;�J)A�ۺ�v
�[�a�yv^�_����U�c[����M�a�U�x�h+ �>D�R�׊�G��q�++K��a�@�������;���W<_��~�P&�N=��7�m8�KI�Il�~�<)��oPz�Q�_�T5�u��׮�:�Yl��Ew��0�ix�)\O���!�C+,����|�s�R�$%�;Knu���;1b�),�#NG\A�A���R�̜����Q{{Zz�g��Gg�iK��X�+�<"/-W�)<�+_,���m�������t�URO��5�K�v,eD/�@)���?A���ޯ"�o��2��];��Tm�Ǔ/x�P�����t�A���*��3�?�o������=�.P�V<��sm`���a��c*��>X�&I7yi<�kt�mnC��r廩�Y��0�����6�����?Ӗ�~�Vܙ����V�%�=���x��ldi�G~-$�Nى���@��[<k�K
q
J�Uʚ�a�"רּ�mb}�R&15�(�
�*T�S����W�o2�Y�B�21z`og�T�G�������/kO�����+���\���0R�N�ҫX	�`�">s=]��{�Ѹ�t~��Q�w4�޷����ۘ���	v\	m�-G�f�خ��rHƊ���㌾D�Ew�۾�w��轢�����%q��Kb*ч19*�5z�����S,mQ��o��l��*QZ'U^��,z�|j
�$�97a���@���?���00`��v����J����w�C!��W8V�������J�+��.��ںǤ�wȺ�"�F�ڄɡ�0�%E���ݷPLjt���_(gI�ܷ���x��v ��P����!v�ıA<y<2,\&���ҶI&�/@�ذ�ҽ������k�FY�xX�>I���;��_�߽{\ ����Y�y#0���o^cѦX��95�os�F\<�����e�w�롋�:��8��ֺdz}D�X��IX6��C�C,�)�1s1g�产���s����(����Q�,`��	C^4�Qb��!Td�11�#\q$p����AgG�_K��('Σ`(^�e�C?�`����Vp��7Ӡh�hR����jyX�Fb���2���J�w�/���~t�*;���AQE�d��F��c�N7ܓc���\�����)��Ql��ȑy�G˂�=xm�u��0����'T�{�t6f�7�o�GJN���R�:8s�}9@.'C)�B��]��&v�&�N0�]�X�	U�~��B����H�y��x���+&ZU��a����f÷�|0أ����՜�g��H�/���fOr7��y�)���F����h�X��ߒF[����F��?=#N�r��&�^��#﯇�c��u�70��r��ﰥ�����?X�l���mp���G�f>���j�-����Y�T$n_�x�s���ѯ�
�J�P�'�=}�[�
��H:�������L�##f�Cu�d��XT1�y��Y@ ٔ����F�@</}���_뇛8r~�Xn���
^�;kU�h;h�ʙ�"��{h1k5�y��G��F!w[m���\�B�l�5q~�g��/�;�2�8��wL.�,SV���:0e����1��:,ܤ���3s�@1O�ś�ì�����>�k6 k��*M[���.�/��<�de�����_�����=]U4N��Tr���+m���r-ǚϑ-��}r����B�\'��/��u�?�$O�KK�|Ǖ)<��	=e��>,B���#��ڟ!q3�p�p-��i��h��wB����T�k�;x�t�M��o��_�Ur������?f�%TiJ���@���n,�P��Yҥ�7�ߖFa_k+嘪�li�?��o�N�r��V=Tʷ�Z�{�q�+�y�p8�ۇԗ��i��[�!��K���k.�yD�	2�S5&H����YP��2�\���)��iϑ��\����f6f�f��b!/B�j�g��)�,�O��K薒ҧ��.�Qu�/X����-3*�'��վ�Al���]\�H���B>I:������
�(�+q��D��
��B�Ck{S��U�D��
 ��(��ʴV=�k?����c%ܩb|cp��V�a���}o��u��P�=v�[�su?�E�2bƜb�g;-E{\��`�fƴ���?�<3�R]�`�c����~����[
L���k4�j�p��qN��YvC�*�(LX��6�h��A��-�łxQ��|�*"R��G�JUk�0 ��+�2�!+�n�U �H^��(ۘ2�����HX���D�����d'���R��>Y܆+�/����bsXnhl�f���`����6�'����AP�a�)84}_���/�l�ExΌ�5���x��I8��.*n�'CyC!.�@Ϲ~�&苼d��*@���?dt�b��� �Y]��/�g	݋鵀��㯨VG�SY�@d���A�?�գ��V1�CƑ�%�8������{~�y5�s���/eNp��GK)�+,��۩%�+֙Y�������-6�X.�ΚY��������c�q�����TWl ��XII�d8�u6�8�7^�t�{�$��y栏!E5��٭N `��?dN�#�Y�~�|.C3>�ɹZ��JT��lN1{��2m�ڐ��s�:~�3���«L��Z-��n����Bc��2�I�m�^�8T2�� +}��Ù����@��Uײ�f�(3�yL��z��q�F.}=&C8� �]� ]-oa�\��"��b��$@��q�E��Q?,�����+Ȃ���%��l��Sܬ�%Rkpq�wg�8gA����ޮO���+kE'Vz昁[�iL�����G��0��ي�&��Dɿ�(����q:�S�I/�r���ܙg|	���#��E�w��{v��N��}��'�te��:WJ�{�Z���uJ��e)�� �|r�F���|eh4�Sq��2m5�T7܂�k�`=��hţ�Jh�K�G�yC��̻թ���D������JvM�Xӿ-�p��DH����˜6��*ɄRh08|9'd���T�i��&2�.g`�o�
�of�ı4������xk#��B�����F�^�#_�4^�;t�3?�}�q�\(sx`9Ll�M^4��n�%�;��1��$#�����g�r�&�������]�񎲀q''&�O���r�S�� �_	i%<�HT9u� B.&���Q�ǨcB��2��>�A��*hG�M��s&�}��LK������r��0P����໧��$z2�� n��q!�����E��1C�=H4Rb�^�^K�B�����k8�����̥d���n�Ya+��:f�Γz��+W�[�l5��S��0���ʵZ��.�y�y�<{X|�*2E�H�5�u$?#�̡'�3�8���ϒ��bFm��bY9�0�J+�
NGE�l��������v�萁'�@��ov�Pi�[�)�g 5���A��xeW�f���@ֽ�fr��H���P���?p{Ps��2)׋Q���a�.�
-ʖЄuf�ksK�ɟ$������uuyd�'ϛW�94��pN��Zpx��h����Z��.d����]���]ʔ3.|���3��p����N�RwS�p�������,�)�t�N�&Q�#�Q�P�����G�wg��ߝ��k�4����l_w�"+k���j���$y8�'�̬�1��g|�H��"�.���ħ����]`�D�5�ז��i�7.�a=����P�Y��2���׏X�+�'q���v6́!�{�`?S	�	I���b(���!���uj�)M��(Ͼa'���A����\W�\�+*����>���Gh �}�V��zl�1I���Z��ٗ�C��v)i���^M,���-���<Ig���H�@f{�h��n��&��N�)�K�?���mum�4����0�\*�����������~�s� )�^w�ޘ�ه�&X�9P"�JFeT��Qy&��v[�����xɐ�8tC���|���,[0F`
&��4Jƪx��C���5�S@����ϙN�١�+*1va#�dA�~&cm,�V~�x�j ��5�����h�>���D���?|��%����������w��W�uA�e&Z���@e��t}�3!�KӺ��ER�2/i��p��i�(ў�z\E��+*���x�����m�n�@
J��5+�A<�����p@v�b��f2W��N�4�Q��%Z�d�C��"D�V��Q�f�������8¬�S�b�CJ���"��sG]3�
��_j�����I�R��3ۍ%�B0d�SVϧc����ď��E�̦;������/W�%��t��Hx�J?j�yvE2)t&�To�y�G.V�X �n�(�.y�^�35v\� &�I�SN�N�0tp���X�r�!Es�{#��+�CN&�������Lr�³����2�	��O�k?r����P I��*�ǧg�ّ:�1��R���'�Ö��fs�0Rl7���ǣ�]��>Iry�8gH�T�@*��(�J�7TJ�o�ْ+˲i2�W?.��	(��!Vܸ�"�אYu��<�R��J������x����
�,}�(�j{�I�q���(��U��o8K�H*�lF&�~��w0��e���r��}��1-��AĚљ[h�B����r�T�ᅎpr���Ӕ�R��I�x���SL�|�kW�y��f�
7y�)���2#ud�|Pf����0ty��J�����9ZS��n�W����L��A07�a��:p{�ܟ�s��@�{mY�9��f:)��	��L�\|�!��R�m����I���./F��N�0ĥ�$���Ɔ�Y6�1P0��"�klS��8`o�z�~:20*�Z��A:���\�O����ו�^��N��0��}2`�CFŝ�|t�Z
Z�9��yt�hN�i|��NT9�h0vX��<�l;2�6&��D�4�� ��1d$y,%K�-,�h��LԠ;�Hs���9�ζ�|�Q��L@J|9
��\Kf�N.tu<���Jy��$�'����J����&�����k^(����;�"�+�ߥ�HIXx�Od�'	2�~<*U�Jex���z>1\�`5C�AY��n> X� ���ð��Kr^-%m�����D�����F,?��Z8����k�~����C�Uծ���I2o�%���nQ��8����,Nw��	� ��`��A@�XT��^�j�YgKw!�!�[���mm[��3���5\@bֈ� ���0u�DFB8���9b�eB��w؜�u�s蒴�EOx)�i�ړ�۪g�����0�N?/�?� ���]���Lv�9��cn�6�{9�Ǌ�>�9���Z�S�1KJ#������Gk�@'��S{Z8��BI��P��������S�Jԝǲ�;Vֶk�r��4����?O�����v�yu�Pwt��D�S/���(�M��޲.�xZ�[W	�f�Q��������Q��(@�Ih8�Pm��1]����1h��ܹS=�����_tr�tJ�b~�uS�("7KiH=�_�`�As�q \[�X�%�J�f�W
yP����-z)B�?HcK*�̒Q�s����
9�T�;�8�:G2�:Ys���O�c�ŝ�
A��Uu	��
'����-,d���n�GT,t0��K����G�!KQ�Ę�xuU��\t4�K,�?�k�T�>TB�B�;�� �>7䲝J"���x������v�Y�[�<�]���.9]=�o}���t�N��4pcg��`�I�����1*�=g?�w�����]���y9ڰR��2��M��&� ��=��V �ʅ�H��ٸ�w �����I�s��y;�:�������r�hW�3�f�+���O�z���C$J2��d��0�i�y�<	3����c�2K��z�p�k]QC�u�e����F3��|x��".�����-��K��q@�����y`RM�^_�ި?)�̜֔e�aCf����\nO^Q�1��}��|x��.%���?o��p�Ѯ��Hq�t������ r�H_kM�x�g�30���^<m��1rw{�KO�eW���C�䁮�������IK�,$��mԹ	0a�dq�ĭ�+�gY�{���y�Y4��ŧKiS��9�ӐH�-Ƭ��rQ�=���o��|���R�	("�J�@�q�
r
�D�3d��$�g��'�'m7�f�q#�?_�H��k�Ke��*1WF�矟�Ӥ�!�R ��4?T��s��E"����&X�.����[���E������|���A�K�w,-�*p�ܶ�V\�߸ڊy3��kZu&(�D�~q��[����Ujk�ҿ?��UqD÷-�د�(�:L�(���fq�kn��V�[-Zg��i�m��{���(һ��e�D��;�?�l6��5��ܱu�O�_�����D�f%�c�2f�51������sA
�͉�#v����l��
Q#���M�ּ����������?{n3u�@�O��!!}ٕ�����) YW��j���c)�)V��6gT�����i�U����!M�d���L�v��""�)%¢�}�����#�Xİ}sAmTY��Խ ��v��tH�k��є"z�ڣo��{�	Հ���0n˗쾐����8��7 @��~�;��I��>�&�h���� �,�¬QW&�}l���2�^ݓ��(���ѣ�%�~�b�]�3��/{<_����dc
=SH�  ��x?vx�%�:c�|�&d�?_�P��$Z^zpD��=��W�N��E5��~�ѯ��.�Qd��6%���8�"tNg���Zg�Wu��.�p^�p�b}�ZE��ޑ��ւ���:��G�6�lc��JyW�)u���췝^�[��u!�Qm_�ΐ{>���t��*2�A�>Bi�Q�;��M�3�����p�u�%xƦ�)�;ʒ ���g%�VB�'���Z_��6��S���R���b�����=G�)]�X�Wd�O8K�!�Ɖ���JGm7�3�{���kW�[�d02zE�2��[O�.8gC��&f��F�e�f)8�&�h��^��_���o��/�?�)�q��cӨN��7�Y����
!Wٶ	y�(c��	Z]�7wP���c���?(��������fZ%�+�뼧?B���xN�@ɯ7��x�� �"���E	�դ�l�d�z�X_G��zIj_�K�Ⱥ|�N`CldC�HP�D��u��$���ذ<�H��C̗��XOõ���P��xn�K�5Ƚ�_��n��Lo�(�g�F��<ׇe��g���S�W��b*�������]��Ȉ͘	w�y�΍������������w�H��RX��M�o��젓]�n6rR_��%�^��M��##�]����A�����F��a����<�K�#�nY��;(T�dE�LS�r�"Y.L�k�aG��9&����Pb�Kwkk \a�Z�.��Q�"��O�jΏ�e���M|�&�G�ݿ���CN�Gz�� !�`L01�kk����2pώ3��z�"?��Ĺ?Y�ÃvPX�i~Ř�Z�T�������Ա�\&�FF��
&�E!*�(R!5~�M��<��]o��ieR-�� ���#��~%�錫Z��3�¤�P	�4��<�+���)�{�+��4A�B�\��)���
��<�Ia�%j1��H
�^E����ŧ��;�%�;8���ա�����I"} pc��j�%V&P���6cCzM�]�1&��^�?�E��h���)6X�]p�_�"�N�]j��w,��@*[��r5u1�����Mҥ�w�;A��D��/�Ž����U)�}1�]S�7Q�f����X��>�+�3]C��W�{�a;�MdY��r��@�E+	MD�/�$�����_�T���T�p�ܝ�e���y+U��Ƞ0>���d	��2��e�ˏ�����+�E�ze�B��aP�g/���K��~���G�/L��}H�h@ElΈ�-��7���󠩞.*p�j5n��72;v��B��|qFH���1h�Uw�������1���d�2GTn��vHZr_ �1?��iRξ�X�~hK	9�pzL��ѩX�t�l�"�{�$�L,ż�װ�E���3N�ߧ�+��
�徆��$e�K�*v���Og̾�`��ʄ���pJ����L2�w{Ï�ky����톃��s��-,���w�+��Ѳ�8pn���l�U�����9�RC�7 4������
F����������ley�IzŰ�����g)8[�)��Z�f�Y�t^�{(�Q;�H���^z9
"�[�Ċ�,,���b��C��$H�@q����H~���({�@N�v�IK3����u��v�]W蔈�fK�l�V��A�}����b3�K��a�l����4 �B�T���"Q��(	<@5\c�g
�l�jRDQ���\4��V�mR���Z܁�a�!.}�o��ם)��?�=�[��(Uf�h	yr��������.��ڃ�lMNE��x���	 M�w�A�E��K~��m���MODr������6�����L�`�ؼB3#��,�����f��0������'��߹跦�0��N���י)̓|��΅��݄����`@��X/���
���9o0��h�{V�:�&���`�t؇3_֫d��IP�����E*�d>�鐾献Z��ʍ����cs����
3���ދ-| ����㞧�50i���a�RhWua4����DE�!_�^�î���%H4����(7����J/2y�(~�3瞌���ZǓ�?A��H�G�"�M�K�n�O����z�$�,������6L|���|��&�LТd�}�<�]�x2�>��4�v N��-,1�:b���Y{�n �"zȵ��Q�L�t[ ��[v��"kZ�����C�~M�!���<pf@������-�v #����OWȽ�����DJ��Gw���K����@�8AC�>μ�����F#C��n���T������+pw��htQ��`0�]�1��h�̞�j���#��֓���ֹ���ꄰ���(���%!����>G��y�p�99�+<`�|?����	'��j���ܶ{z� <�I�a<�.�����pC�!v;���f�ROS ����nȂ�?�S�b#��$h6p:!,>��L0ۍC�#VkvKj7D���ɛ����*�����Mx���z��9E>�!�1��#W,��p�B3���?�V'�H�_TwL�i�8�>�O^ @΃m2��:ۏ�"�B�r@�����Z���t[ʬ�z��O.�:�}e֞W�O�9��+#��J���v4�Z��ީ��H�L�TM�`��DQ����(��a��(=�3�PbO���= #-��^8�&)��d��#�Ql�D�*�(>a��
��B�a�Yٕ�{�� &�����w��i}u�k�&(�R1cL#ڬ���Q�(V�̞
<~
�41\#2&���E�՜�e�R4�N:����Ӯ_-�+�7�%���29׻$S�/��;YWG��do0>@��c�WíA2������EV�X#f�ߊ����_s��r]&��#kP��R����_j8x�f($5�1�ښ�!�dU�C�g��u��QƺH����Of�
e&+Fw1y���y:�p����(r�7W�{jY>E:����#y�\�`�ث߇�u��~�]8e��'L׭�z�{
�����hB<��~����%��l+
]A��q÷om��=���ԉ��`�����<�z��t�B�%]��\�<�}?��������.챗Z�-w�'o0u�M�hio�5���6�AƋ�	��Y-��W�y,���wD����+�����v��w�pPP��I�o�Y�`�x�*��������/����O"�/�JQ\����T�4}L2A��Qճq�.��m=�z���=y�Kx`U(_!I��JQ��#�7�T8S#ɌƼ[BS���j�N�E�CQ��o�"l������^��ImJ�}R�	�☜Ģ����@)ل+͠�[ڨҴ�H4GFD��$/c�ƈ�_��
�6�y�o��nag)�4a/�v8J�ıpnC�g���L�y��,~���O!a8F���悋m�L�V%+J��;���
;�3[,�%�D+��/����I�-���d�}�"|���Y�_K�UR�D�x:mK�������j���y���9t"��P��) d�a���LP�v�c�2��1�yV`Q�}������Wg�`��[���zǗH�"ON��]��y���A0`���k+5=�>8Q�>�
S�����(��E! �	+cl�ree=�I�v2Sh�����<MSZ�.~v�U����ר�W}����Փ����%<hq�x.���2��{^�����1T�>�ST酱k��Ro^��4+ڶx#v"����0�r�o�L���"��h��`8��p oa��~T���jZ-���OA|�]D���v�@���t�W����ɵ��� F�̨�fR������V�C�G�m�{��[�qE#q!�lUI�$O?��}�B����8�&9��f�����ҳ@8J1����lW�0zjr�D�d��QU=�3k�����6-iG��.{�x'$7�/{̖x�&��SNy>h"�p��| ��4<�S�"@P/����YIp��q5�:EI�Q���� u�Z9Y��(�M@e#�$V`������� n��%�����tT�8�Å����C������ՠ��d��"Il5/[�:���},<�]��3��#n{f-Ζ��o(h+�2�OB��aU�z��7̤�#r��A��)����Zuܕc��"�� �A��Q�����
/�u������:�����)@�K?\��-��X`������k�yУ�3�+�͎}i�Y3��g2�I�{�֭Jx��p6�)��6/�15���(��0i�%�<�>������m�keDy�O���FnW~��p�۞�C�d8�&� �n$Gp�ɼ�E�Nc����O�^�>�������R�	"< �~{:���dv�6't��}~�I�%ɣ�E�xi-����#��uAw�����ڙ�N�FF2�����N��@`9�}�3
��gW'��X��P��m�6H�u���-�K�&a��ם�j�b���� �Xv�YH��� �Ǖ� u$��?�����=D1�ƦOFf�#�z�kD��1���QJ@Zj�J�� 6t�۝��K2b�I�GW� �P
d#���m�-p�{ �DG�!�?�>�g�����K'�)�۵=ehQ�`3{,R�����c�U��@O~A
�ŵ���\k�86�8�
yߎ/�.8W�Tܕ�y�-O؀oE�Y�3����%����;������r����=뾥@�X�@Ź�V����{&b�T?>����5?��"I+����)9AmI�Kc����w/*OJ�#��/��E�*733��d-�fv1��S��(�J��m0����vv�>e�h��"��c�[,�֥)!D�q�����{�owh���^dw;���i��	>�6�$��o`��'쟎BCSݤ��]{���l�al��Rq"������7;�8c�l�|��u�W$�g5����ZҸ���@�N��b���xܽ�qmy�Zg|+���q����iw��Xzt^U@���)��`�����Cr��s��#��U�T)����<�9a��u���]P�r��"�����M�m�rT�@�GRu�sT�n,f@W���*��E�A����^t/v�O�0H�t�TÓ�k�v�s�6࢓�"���2�'B~�,_���b�&5~���=��5��Ml~Ж�1F[�:�w?�[lW�|i�j���P�t�x�oqԚ�� 4]pEH��M	���C�E�k��-�W4"
��d�|o�v��oP��NP#�5pM��z*6%��C�x��$��6�2k�Hp�0E#�gh0S�u[}c � Y6�]YB��P�����)��h<��0</�<Xw��9�-�;4�a�ux��M���2�wig�F����>ؼ:�S7��CH����>�,N&^]z\*����WֆR��Q��?IS5F]ݠ�&a^!�k���.��ge�5��c�&[�j�4g���s�>�e%�e�a(�f���I��d����%��Ƭ(����!
����|�245���֮H��&����[J=�qwr1�\z��q�.�Ȅ���)r��`�§�9�g�W9P]a�6�ԃ�uCXU��[��g'x|17ֻM�c�x��G�:���/��\O�$�b9m��F9���\vq����]��n�}h��K2���#��:�$\����;�rD��)�wa;4��2�,[���`�cs����Wb���#��>	u^-�Fc�X ��DwT*4w��4`��U��I���eYM9%8}�W�T�U����� �rfDߺ���ͤ���J��-w���Ab�ܿ�;��|��z=�4�����.A�Nx3�8V��l\�>�T�~gQ�'������i��Hظ��Q�e�����ch�ǆ�2�E���F�����d���t��U�;8��p�/������	�Ŕ��7?�[-�x��A�ӫ��5+�ʑ��/��P!wy��Q���.�"N�����V�[�?�&�46���Z`��d:�+M��aP:x4����<jM�*��.�@���ʑ9'zR�焵�R����l)�8-��MHY(�����~d$�n5���B��;� ��3�IAP�z�c��r6s�1�m��]}C�#��o5�z����㥞�E7x[(t6������(�{�_��E�΄V��M���j���g�y`E�t��U�\����/�0�铵
 �#Qf�M�$X!�{:�!,��#<[	\)��Ύ[ǝ&�G�!�+N�߯#����'�|�Т����<�j�L�Adp�����:�aG���GQU��s��V�ל� �1=Ha3fE	Ds�l���'�1V�j��`	:t��1���Ā1h*t�d��kD���Ƣ�"8H?�6����nR��'Z0��85o2(�q�/�z�-N�K�M:��)�w�`K]n�M4Y����z[��STp,V,"��5�P�a��l�U��b��&�fJQޭD"�-���jzlў?�r��gg�Ŵ^V��rǶVg��W	�G���alo,l�?YQe��p�qq9�D/��Zj���<D��h��6췰�^�E4��Ճn[le׬3�����.�;N���Q�:	]�}@y`U;O���(�;JgbX��Ku���$���i���u�U<WK����塉H��Ӹfq�0��I���Ŗݔ~�<�ӱ
�����B�X#�TG1������@���!��sm2�"~��V^ci�e��*��q�y{�7=6�y�[�AU[M��wJ>���K��6�cG��]\�S���P6
��bZ�Ce&�#�Y�$�D�i�U�Zvz�ט�� ����0��`��Z�N^��	�����H�c~�q�1���
��dPx� tj�S��m��]��i>��n�A�K����c��b~\!Z)�<9�sn�>�����85c�Ɯh:����\��'��5���~��P�^�De����MQ��dN�O�������Q�mU��s�= �Rw���6��\�ZO:>a�˷ރ`�y�E�qjIǗ8� ��_����d�#��rw��4f��8I��`��[�=����W�Dm#��g�&Wa�aI���K8x�{{�BNvh�l� �L&&+oS���k-4��,UA�3�ҪT���_��뚳�u*����P�Ky6vP�q9��-�� T�\~׬g�N�/q�5���l��l-4��q�]vc�R�P+�֬}U�X�˔0$ü5Tq�E���H�,7�f<Z�V,�Giܕ-����q��?�N V�p��D�v��o����Ȃkz�0�yH8��]7?�/p_нu%HѠ6H/cρ<L�=4o3��_\�p�1�!N�B�M��d��'�q�����������jo�(aKe�0�ԣ����4ٕ�����1�QoR2�D���{����tBmf4���G�J�2X/�b�S�^���<�
&���9�&��0=9�/Z���(�v��?�M�ّ�%�E#C
p>�[x��>����r��o*u:B_�=�+ȇ�!o��L5>�wvw��2�b�>{�e�����٢<�Ɨ�A��oA��|�� ��ݕ�����8�yU��@�έ�E޷�~� �j� ���j�*��c��%��-��V9#[K�{#�8'm��&iC4�>߫��[��
������m��^�'��l�Xه�{�m��ǟ�V��E�L��i�J�0%���V��{�Wl��{�����ձ�<W����KR��?�wa؈�?u~{}��s��B�y�� AK�"������F���p<J��F�Q�Ûe��>Pd����A3S�%m��>g0�<�Óh&���A:�;��ElA���1�˓�����\���x�K��;��Hⶺ�ǁ\~�����~4������EOv�	�1�[ʠoúX�Z��"?�_,�x��J��@���ҋ䱞��Wϗr����!��U�|[Y~�:=Px�@�Νn��QZ��s��kc6W z�����_�P7Q���Du��e�y�ZP�Sv�.�4�'��v����"5c@���9�Qٚ3$k7�(#��v�"n�,L�a����Q$Zc���M"Z����9��fT�H�8��L��E�7RZ��u|Q�j�T����X�~{W�Ri��e�#z�ܗ'�[2 s�>���z�̉��2��.�Z����87p�}��'B��Np�,�����O�(��>ƶ�Cٟ�A�LV�&���ίӉ�X�E��l'�Fs����vK���X��]�K�#xF��F��jV3ƾ�	���O���o$�����Uv��Qs��żNos�@�+�4{+���U6��u�Ҧ�&pؗ�n�cN�2^�'����'y̗M�"��G�gɦr��I0U1���4�*%�?��0k��)���f��xn�Q\�O�B�*f�>#���%3t��ު����$J	VE6��%l�}�4�X�s @.�Cl�$�v�X��'�Ib�p��b'Ɗ�6W[���2��Nf��0m�"�Udn}�N��_���D��z���!ī��b��#��E��o�[	y�!::���ڲI���y�Ԕis�5c���C�����NG�P�Բ!X�;f�k�G����\U�5oj�1�YS�(,!�k�����#G(�b�H�bEU�̾�e9��)�j�����?.O(R�{ug��n�:P�=%	��NT�v��e�l�&N�~jȆ�qo��E[KyiN���'  ��aU�O�L�)k����b�缥h��DOs�&�{�Z�.�:v*�63���$ؖ\���P�B�5=��+P2'�A����I���DF���� _Yì�	9����#�h��y�a������>�:w�#�E7�+�+�F���\�����l��:4JG*%
zү���}@�I�"��uVŞ%R/=<M�F츽.
�|]#�ؼL�zX��9DIWLL/����:9wݥ�?���;����x��U��_S�b������o�r��<�3u�
*��xR���&z��=��ܲ��ī>��8�W�p,*��N󪈰^M�{W��L�6��o��-�O�v����P2�o�a�q`@|�BDm#Z��r���|x��ȟY���oF3�9>\��n�0��j�ٗ�������"��z��,6��i��ŗg�f��.�,�?��3I6M�ةF+4 �1jM�L
ZG��x3�w����2)�O��M6�꓀<x�7$/zGޔ���2��x%���ʅ�׋�;w�w��6Y3L���� �]	и��!D�3j����ӈ�a��Έ1=f����)fO��p ���u:�mrM������~݋����%w�W7��­�+ƭ_���M�C�a�woB�M��eU�B�@��Wt��LD�Qs�������褖"n�I�D���d*^��P�-�G�JoV^��N���U��}h�bnBG�4|�@�����( ��t����ۄA<���fş�Jf,�������B/�UkB)�������No�3G{�!%a��a���!B`��8fb�]��6�ê�뼎D���;!�D ��uk��ake�;���E.*�5h?%��&]3
"�4��ƪ=��g��ٍ�$E-˵����/�T5��@e�}��o���.��ςd�-25�'�t�x���1�����H1�cY����}���@^Q�����?�Tn�����3�/Lv�=η�8�����MR��8�*j�k�;T�<�n�i\x�Q��3j�^ꯢ�C�	�鄮 ���;�>.<�@ǵ]yg�g�;��C3}�c!T��v��Ic+K�)	d(�8r@�~�c[�>\g_eiі���K�=}ϐ�Q�Z �.>�y��}:\�=�҆ӽ��׉�E���p!P �ƻ/��O>~�9�_�IAw4��Վ�9U����~�+�{v��1{ΊC��h��&�.����K�i�#A�`��>��f�Y�Ղ��G��{��FV��{������8?�	ǁ�Y^�3�}�^���I�y��@�ۈra\�^N)�Zmei��/����z�d"������ex�R�G��oT�,���w�9v��h
d��M� N,�����Ȑ,<��9�0��ƿr�U���yZ5��6����A���G�>��\��Yh�W�%�l\)a����sRНW�4Vz����л�`��VCbn�`+xn;9}*C��p���;����7�{�"��g��<�oO�����Nui�������S�\*���7�.8�|x^��j!���v�Ѥ����N6 ��ǋ�q�gO��-r� ��Or�bS�'�W�?�O���,�����c�K��&[]�I)c2���8�7��;9ܶ/��;�C���>ʿ�8G�!n�D�l�x�ix�p���L�N��m
� CN��f�e��ےm؂���}*��~��! ~)��/�.���K��&��,Dm�*;�H���0��B���{��ebbN<{����$J�ʴ�*�V0O�Օ�J֮�1ap�^��ya�븸/��}����KoĪ����`�'x��s�9-��iQt��u]��L�0��t.�YX?>��dM���zcd�.�v��d��Zx՗����@[2��Ji����JTB2ٜ 	T�M�U��Q'7��Ze�I���{4�B��2�|�q�4y�ܣdD,��ҹnK�S��q�t�ne��Ƙ�?�L����� j{�I���CΒ���gէMZ.���ݑ�^�g��_`��)���Y��y`�1��9lvV��Ć+̺� ��曇�  ��t��p�Y�U{W������Ԇp���]�;��YZ)D;�Z]�S�..&�1+"�>D�7>G=�������f�s`�K�I�Yh�t��=S\�Q�&;�\�w������!Lc(��/� ?~�	� D�:І���A��	���J�:]��^�ӎ׊uճtu��^W��y���j!�~��*�����`S��h;16(3��`B=�|�QEwRu���ܛ�O��B�c���&x�~5ȋ�!c��j�<�Ǽ�>f�����XX;����6[�3���1��LAQT��Yٯ����7$�<�!��[��T6;s�����M��oJs
��Æz�ښ�0�s�L�����ǽ}������Y�dW/�/C���]Xo�ɦX '	�A6;A;w���^�@S�ɥ�j�z�]
����m'Y�N<� �շ/��a�;Fy.|�����g��2c�r`�1�I���V/ RE���\��yK�����Z,O��"�1
�
@��?�P�[�b��a�ѣ>5���$:�6���%�f�t9����RC�J�7��V�pG���-뢝�z���Lդs�����]X��P'��B��r�y�O&�L}d���[�FYV���E���wJ!��~q��D&��.K���zH����Ȇ�O����^c��:��eQ����4�p�d��	P��ܦ�ko�ߖb~�2^���mUy�*Ql���8�H�oZ$IB�$���0������yz�`�5��u�+]�A
���e��k{o	/u���ye9::��RD�K�K��]�ў��y�h���{9�/R���a�>�ퟦ��$�=��h2��:��s��i#�������уR�vj{��\��ɀr.���tD��O���OH�+:6�[!ly��,���.+PE�y��/�B/���W���D��d���uaf�	�o�::�pi���v�Z��nM�K��IC��%+3(�8o�ޖř�����V%���z0�7~{�?&;/}r��+{cb΍ڃ����� B���	�L���i�*�}�_�v��:ö�
$���
�:"y��NkQ�s��b{�e>5$��;�=G����H�<dM�ŉ�[�w����\��x��3�`�
2�H��u�vv,ݯ*E�vp���s��>r������ٱ��ӢⳆD��l+@y�AY-6�k��r0� �M��G\nY/M�_���/^QͳO��?�:1Yk&E�s�xAL�Q�>�:����T!�\܂���yy���Q���%� ��x���!���"��s1����Pm��!\��"M����1t�+��������^~1�qôU��`��2
�S�o��Ɓ�#]�u�_�>Ѥ�bB>�T�:a�U6�o�T+6��uthG!VA��G)���$�҆^m�{���<g�)�0[�ҍ�㥁G��9��/T�æ~�l���~ן�8W���k��� Dd���X+:�^��JW�Y9�ox����r�z'.�������� 
Ovmf�����,/K��]��fbH��zhϱ�D������Rr84<xb�����ܑ@,��xZ��YD����|q1��c�Xx�t<W�٥�A3!h*|��B\���u�#dB,e_f�-��PA��eB�*�'HШr�_�|B��!�L��w�<�tO�%�-�o2�J���n,7\c���\yν{��@]�XQ?6N]������W�FG\�>l�#�f���2o��q���YU�Y�9��u��^�WCF�8�2�t\���S�<�Y$(3�9�}�Wx'A�$��������G��8Aqަ���AbR�C>i��>'��K/�uxK]>���D�!�I��l��P��8�a�1i��/LҜ
�V3��Y�mAԶj�H�P�._F�铂9�˱ч������i�X�#�K&ߟ�y��R���������_���'��~�K�i���j_ G��Ftʋ���9Q����Ӝ�ԮK,�f����ǘZ06�-v��V�U<��C��/틣����O��Xc��0Z�_̌N)c�*b(���+A]!�ݬY��n�5&p�Q������卐`*{t�qeg$ʦ�����归��eR�q̹?)�ή�d?*L̛�}r�֓8����(�����s�Q�i�rr�)�!l�M`{?^��d��~�z�[�_�m���U�N�I��+���l��//����[�������U��e��G����9� ~�^�&�$Ӭ��$>�Kܬe�������*��-k_����n~��
��ƹ��.g=>�!$��ՙCa?<ݠWU�!�q|�w24=�@�W�a�Y��'w`k���>/o�Y�	�]q��tX+�!P,̮Oʒ��U� ��~��7&/VI�YK�-�7��\l������be�yE6@|+�Q���+Lq��*�\!���#B�Ʀ��} ����rW>��Q�In�8��,��g��]Ѯcڕ4۠�az.a�U�Ȥb���k1��A��;���=>Dy`�\F��˻�$�0��
��0⢱ ��	���g�ĭẋ����~\��aHr�����7� �x��bs�9�B������0�"�)�_떊��Rr�:�+ߨ�Y��n�v!�K���G�"m���!�
��2��ۧǂ�V@��4{��5�?֩j#rh��cu��7)Ө*�yꅹ�?�0;l� Y��j#ob��%ʁ������0|z��$+�:��'`�ݗ\)�h�pA�����U����������l��t3�u����*�ւ,Y6&�Cr�J;����V~�8[P��1'"��Q��*����G�S�5gݢ�����@Y�hQ1�
���Ŀ\<	\���,o9��Q�Z�s�D,��,��R1d��/c�&�̼7 @Ce1�J�^�b���ߌ��&��P�������3䠮T]z�e��W�9 V�ղ�d���P�v�IC�#Z�:L]�a���7G���ݎ����~[N|a6�:����W�,�Sʙx�I�S��7�B�/Z�=iv`͵h�B*0whNl=ק0_��C0"������}�G��9a�9�9`����G���!���kJ��B��ք���^�}�:�Ë��f��rL�_��� ��c��F�	����(5�X�%���6�ˣzݷ����nt鑰 ���=��s�y�H��-�6-�Ⱦ�yߥ_NC�髥�>�`
n ��v@&\���HS�Ψ��v�^��\����MM��9쇙3	1�w���Y@[�}��>��^�W{�?%�%�;�4�iL�~}S:G2�p�sƾ�*��P溺M>�q^%�_�0S�m.�H6�B.;����7���}�YƲ)��Y*���콧$� ����6�-���ܫd�M��,�fdq�_��?�_�FIi�G��LjG�Ƌ�r� ��$���M�5n���P�Q䚛}kڥ�N�Q�*.Ux�ÜZBdKU�y��"�3J��]fP�K`�� ����+������:��6!���/����5�6'�S9��i
������q)qR�ܕ��H�D^�.�X����%�gu��s&h�x( eBް�1�� ߙ6���P[��U�<`Uʵ�2�L���
�ZO�����N�*�������,���0��}F�9�e�Y�D���5k�X�� $~���1�?�Kʨ��F���Z9�w8��q`�����~����<�MC�@""�!�ʠԎ9� В�L��"W�@.M���Q�q\�$���;����e�������6�B��,8y�\c��w���4�6�v���]$��
$g<�̶np:��2�v^���b�K�ih;� Q�dr�:M�����+��ҿ��#j�b|J�j��k�DƋ��cZR�S�j8��0���>�,�ulQ���o���*f-�/�ٞ U- g4��r��Rw�﩯���B���sΆ߼�gʋr��BF�j �s���1��f���.N�ʑ�Be�w���������1/ ���T;W�M�������ZɒFH��߆�D�Et�	�B,�ss{��3�M��K� �us��a�ȏ+�F�M_�p�7�.�>��x�G���}��$R�i~ἵ�ҝo���	Qä�7_�w}a�~�{ <`����<��]�*�J`p���;P�+�����Q�3af/���z�3��Tʼ�E����ߍV��n��Ē�ɦ�ړ��?~�Ս���jӍ��ɲeRxt��&�����A����4R�4Ϙ�f��:-�4),�+O:"eof�Ǧúv����Zk+�!��B)�j>�ԏ�KO
�����e.����$�
b�M�JPJU�9XWN����DB�o[�����~�~�	���=�I�f
Q�h�KM����J�Bm�jF��.���t0��~R�ĝH�N�C��W�/��E+mY�5���}�TB�,\��#�^1����l8�%���q���v�FҌ̠ڐ= �PJ���O���{�U�
R��j2Q�K8HЋiO�W����	�V�i>O0�y�bb!���V��y�������S7[h6�t6�B`����PLg~�hj����qy8�S��0�Z�_�Jwg%]{�F��{e"|�R6*�\��!B�9���Yi�J�;e�lb��R<�E=��?'��Z�	u�}@�Z�捞�F��i��%��B�G�k���/���T�1��B�����۩��[~yy44�.d���"����˳���d�R��LTH�k�f��ᬤ����B4!������y�>�e��"� c\���z��f/���3�4�j�jhj�L`��<�x�r��#���%q��TkE�[�Ϩ�����c�$�Š
C�:\�de��^1��D0�o�]����N_,�m(=d�I	c��@�:������x�A�C�G��
����.���=�~V�YЀeЃз�Ϯ���?�<8ABB����!U3�f'��-�@.T�7�;���c^�j���	��׃)�2�u�T�9�݃�RLM)2M�w�!=b�w\dՋ�z�qd��&$�����V��n���BfBa?��8�keh��V�Y�:��w�*�>j;�B�o���� q���Ҁ��|�����a�VE��N��	���Ռ{�36���k^�X`H�n������<S�d�cZ�	K�:0�Tγu����'=_�=��������W�ނ����G�֩0#�6z�ɗjQ��
�uC/j�����<�xN��K���23qx�w�1#�ɍ��"?a�V�1���s
�����W�jDg��vΖvD��S��z{�8bi$��������>0F?w8bGY�]��&C�s�j�0��z]��[)��-B:��'l�*c�c6>J��5�
�!���9{���>Ġq��29M���y����q�HQ����m+p�醌LͼD�M�>>�^�g}�1��l_�No��A]�#.���'�� ?B�6��.��ӷ����a�?�jt�S�� ������}��Rh��c���O�ۦ(q�'�[�;W�a��M갔���-?�ɚ�WmM]��U@�ڏuT�K�S�0���e�T;�cX�F�ع���K�R���]��d�:i��U���1��J4�P���68�5|�T���+>�j��
7��?�&_�/JAK/B�ږY^�P��ɡ��X��jF���A^�і�w��Q�-Y�U��m�����m�x�=q�U�8g�5ĭ�Ӈ6E��q����#��[�}a�_�ȅ�[Ni�l{V�O�q�4"�y-q~t�	��xڸw�%�9ڝdiy���"��-ó��%��F���[~���&�eAe‡/�j��.,�yPa�O�+V�g����m�J��S��5�bd�!&��r�_6��)�`�X�T���Hy����i �Iw Z�c��F�l��A��Gg t,Nš�@����.��Gn��Ef��ڷT)�kL$%u�K��Ѿ�e~� (�=���2��d�Mא�i�:,խ����#^�*B�pwT /�f̓�>KQ�f�����@�5msJ)�����_���R0T����E�E��"Xۣ��H���и����2{���:��;�c�;�3K�u¹+�ds����.I4�?�� �3�V��X>I^,�H}��My�םQCl<'	S��V�,�l��&�xS>�i���10U����MP�(T���)r���t�V̆*r�*�7�����^���u�X�b�����+|�?�F�
(�-�I<j\�d���'	��>y�;����*g�CJ�!����2�Ŷ|�\��t
��H+���s�-h�������V���H��?0C����ewY��Z��:��C qo.Q\U*o�%�9s0�������49e;{(��ݤ�YfvR�1�#��,�䳂3Y�(���r�UI��y�����T#��b8��H"؉���|�Ρ~�q���F��^��.�V�)Ej��i�V/�tM��ǎI+�[�;�c} �P1�*y�B����Ó샏��;��	����9�M�h�r��p̠.M���xl�|�j,ˍ��R%��r+C�_H��sY�~3fR�zT!\ln�Z��T ����^��q��5�K��\��Z׆,���F�o;�u��b�JԳc4�P�����4\��h��]��i(��|��!�%�1�S%4�G߶]򼤬h%M�\�n"����]��x ���:�6��+	s<���c�#u9��3 }l�Z=p^���r��H���W��?��6c3�L �|i�FR2U��L���t�G�v�<�2jvy$�>�D�a�b��>��o���g��p�����]}h�*��JLO�{��a�.l����1}̗b�wh-\�K�-1�q�����Π��΅���}ݥ�Lҥ��f.=`>���\hZ��M-B�q�V,c���A��-H��)�"u��i��-rb��e;�O���C6�g����E1ɱ_�ޏoX�J��	+�:�J��a�w<G��%g���{R\bFՙ�^Xpg��k��ܒ�ʦ/�e�xQ��Y@�s��� �ë�[IJ�#��8���
0�-8�5dzgw6a"�6z�"/���Ӿ��|f���@t�RH���-�b|��A���(�%�6������w�Z=��A��K2F�#�6(�����E�	B�7��0�l��#t?���G6WQG���n\Sڑ�)G<�3^�P}+.�5c���)]���]�%�zq��#־��w�)���%��Ly���X���I=�L��)�)�,. ��R=� �P�a�(���G�E)i(t��|-}h�jF�U`��e�5A����[l�fj 鋈�$z�+�f�mA1��C�B~�D�ǩ#�`��|!)U�R����'*�ME�W&�S���G��L�8�o���N�c6� �Jvd��	�QJ'��v���;6�2Cj���ӺE��Gҵ�R#��8Z�<T���X�,���Bd)\�.�otue�o�@��&��>�~Y�9�!#��Z�J�!4����҈ �H�&'SW$+�+R�o9�/�]�{�ʬ7�(���] �g�<U�g+���0��組Gq��\r&��wɩ�.���j���0;�X����Y�����?�m�-�
�n���dg��c	#Ȇ�D�U��h4���Y�A��!���I��
H��5��O]f+x>��}Gb6T��x��h��sɷ���}�C��׍��t�3<jȪ��j�f�Ƭ���^l&!�-�f�x7�L������R�K���@��XP�,D+$�#��"?p��t�B�F.!��b8����+��!Ֆ�[�#����y�$�i<k��<K����X,�i����Eզ ���.�]��N����I;۴�b�S��O����
p��HY��0������s��g���]�q�P�h[�<w����GM�E���E�{a�"������C��ٳJ!{��ϱ�,��Η�'��>x���s^�Ǵ����qcV�e���ai������I��'���rRRb|�B���hנ<*�4�6�c{t����uI"��r툚F�G}o���̓��?�(��*����5SR���W�m����BW蝯�!gu�7a�B�Ak�\�{ѓ�ѫ��}|I!��z:N6A�xHmJ�nۯ��LIx�)� F�]��«e�V5v)G�=剛` Ԏ~-�CGS�6�h�1#�ݒx��"�>f'Ndeb6^�W�8���=Շ�ᑧ��)��þ��
��z{��*�/���P��FN�\������'�^g� �?]4ƭ��kGe���u���*����:fBϡ��'-�+eԔ�ٳA���l�8�Ô1����Z���=��i�3Z���§.|p�as0��޸��{Au�e�v�?�˃�T#��D�Q� qՄ��Ӊ���1-��H��CV�`���
;A�3*����hE.����t$\�8"bS�p
��ߕ������e�����y�Qu���I��bz8)GE�t8=`S�W]�����N�dZ(j҂�/�KL&��[�N� ����B�$�Ɇ��X|�<,�\��\Yݔ87�O2߁}Y@쒍.{��`�3#	Ϥ�a}���*qY.�KA<�Y�uI��EY(G\��~����p�UuA ����������U�V)�R�����h� ���қ�M:s����}�qB��d�]������m����Н:_��j:7����d�^�*�On ���²��fL]Ϟ��x����Ϧ��>٘9���&Ӕ��$g�P��	ddF(z޹�sI���\Mz	�7�A���+^�Щ�'Ӎ�&��X�ż_�y!HO���I1cŶ�8(2��Y�I���5���uh���I%V�`0�*�]o��E�nuWm�/%>^���	 T�.K*y�zwV8$o���=�-9�9�f�$�μ�}��$ޅ��U?s�^��������\yI�]}YE�jn�.�C�����iǇz4RN�I�^Sd�-N��xU�Ag�rA]�Ԣ>�рfK���85��E�x��NoLJ/�q('�ˈx�i��L�;�$��z�0�wo%�O��2K��#<GzNn�L���\p���=�<���bgb�91���?�It��QV��U +��E�X�p��̲�1�S���rEP.S�m�.殙Ǧ>./X-�\�/#�g�f�0>�~��Ũ���N�~~��!�@���X�H�ݣ�A����&�`�E^�ČA�P��ޛ��7��k\�
<����"�e�w�G,]
�w?�.�����{mkE݅�e2N�Rw���0eU��z�x��y�W3	���%ns��-��b����^a~gs�������ש�종.�D�dݕ.?��"���s�N�����÷f��HU֋�まO]���>���_]?�KvG�g�k�e��;տ���s��P�1�$�J��s�d�1��f؜��LhB�ݒ�X�5,w��{ޅ_V�wߣOOSQ�1�����,�Ϸq ~�PȘG�\�g8��+�}sUB��_��9H���j���4���fE�#d�dU�eH�������`$�aV�|�|�-��,����OPq�un����x��U�b@,�t�~Ao��͉����\'8��Scx'#УT�_��SY���@����0+�O=4��4��(��B~��(���^�0{��U\W��$I����6#!���1�S+�'M=���s�f8��f�!Φ�'���SNy���'��V�*j�"h���&~W�w��\��7DZ����Kpy�[�,_���q���)�b�/6=�{�Ak]u�c���^"�#@��?L[����e�ǆ0�����{#HeQ��D�/��sB��mV�K�?�#�Q��tD�KKiM$w�&�]܆�c��%9C��00�wK���ӵ��?m�}��=s�h�H`�JZn����T�ux����|YpTW��}�Hc?��E�q��h�w�B��}�͂����7@��q���Ε�yQ�[R�5�EZ��C�q�fY� ����y̮�>�z�^�j��^U	+b�le�>�0�k��ο��oy��y�O���tj;��s/1 ��Ҷ|0Y:C�̹��x�>w���M�:���V�~#�H��݃�r�9�o��w�%��α~P|�+�cE��C5��,�(�xJ�(�|gV����J�=�����zs��F��N������C���R�+$uz�H���Z`�E��}C�-&2S�?��\��*p��� Ȥj|��-�2/7#��X-D��'�O���umb�h�+���=���b.��c�o�����z��s0���W4Xz>K�N�4)Ւ+\�O���^+L�6&ra2�bMО�ȟK�v�~�%�	%#�]K��ϩ�F��#�L[�dS�{z�f��|h 7��
�JV"�����m�f�	���0uZ���$þSç�7�{�R<��$�{ߨ���4����Yu�+���'�M�����v+/{��"��K]�&4z�x�d^�~઀� 1
�{��;�y�� Ejg��4l�N�V�Ҹ{RҰ�[	�@�>��yQ(nDe}w���5�UDDq=�ij_3󝡻���ǜ�C.�W�5B&�B��c(��d�~*��%>~Dv�GD�ӊI0}9w�V8�},)Ųc��ö��~e�Tp�%t�ʑōH�m�|ۢ|�L���2kMhF��?c?t_P�>a���?فȥ����|�r��R~yU�2�����+;A�dY���I�#��o1W21��PI<5T�82�Ջ�_�:TRޥc���I�!]�>�Ƕ��YrixE��l	u*��ΐ	u��)�ɖ����?"i���~o�㴏/��Z�,�f%�$��KoT��|ǫ�j`M<�7`_X@f5�<�bePp�����KXW�4/ωȭ2;�A<����I�L���%Q��_�W��j }7��3�"����Rl�'\��@��I8�Ѡ���N��M`Toq-)pև�䃑������Dia�w(�����j+��!հHu�/�6-�%�7Kc�!&~�C����o�L�K	_�H����-���
Ho]]Q���[~�����*"(�t��� �;�#qx���AL�%�=��m#`Q��[��$���0*���cN�� ��i�7䓱T{�0����%lC�v�Q����`Hsoڤ�6�F�5L����C����}���[�Z-5d��N4�i�ƈ�`��	�3,$7k]�v��}�b]`Ƕ�]���֦��cb��;������e�`4zTDfg�ޓcc�.����j*ǴB��6=���V^��Ua�>����Dǧ�����6��Zf�ܹ���ݑ�x��\��˱#!�&��魋�%�1�M��k!�H���ٳ�ژ�BOh��n��Y�kqeJ�ߗ
d�+D���fK���Z�e&�WO�M������|�'�<f�'::��Kٖ��3V�XH �؅`6]��7C�I��cW$d����ooۮ�wɲ����8���>E�/Z(R�ָ��#=�ױ_� �9�l"�k�,/Pԉ�����6���@�����J:�!��5,���M8����ɾ��1}�7�wM
�;�YT]��(ʘ�����$5Uk�Fx=��Y�a�p��/Q�z�b��~��uP���}8]YkhK�7�A2��zۻ�yI&�D��(M�%�`6qaCؒIȹ�������!>����(��봀��t��ڋ����l�=1$iW;���i��F�E��Q�$~�;U��"���%�Q�\�ɐ��ƙ�"�z����������.F5�d�댁ҟ�3<��Z��8��6 6�����5��)�' X��������!#��&j�u�D�����*M�}��W_{{�Z�O�B��T[̖c�ѵ`n��9՞J
�K�!��ekE4MQ��j Ξ<a�4{��>���P�恩�i���V�b�Ă'��B�w:�v|�=�Y.4����r�DD�ͧ�v�]R��'���'���_3�hg�T�z6�6hͤ�O��*���<2�>ꎖ��6h\�F�@r���ebh �q]�?IF����"1���b}{�-WoG���B2h�	�����wD�.M�ܫB��ǌּ�Im?Ue�s!+�iH��?�oZ+�84בtk�~� ��������p0�4Z�E��2t��]���Ӕ�+����
�8m*a�?�p�1`��uV���*���4�`%d_�3c�='�#yfw�'�(u�6g�k+H?�0���k�9�h��Kv�Cv���ǩ�࢕�̥��pҗ�h<?�s�o`��WZ��T��][\g�G�vF�ꥬ���GZ���!�Gٞ)#i�S??�I�z��#��]�Z����Q�]�+]au��bĂ����<�}�Q�i)/v�i<��"���?Wm0�^�ᥳ  (;49K� 6[h3/���U�XA�\+av去>``���$�Y7�/Q�����XP/!\���a�p�=XG��':wQ?�GvՎ�kǗ��J� �k��6/�䦹�8I/�qױ�<��򄡨=�����i����S� �Fn��U��M��_�w����Wʇ�����ǓB�_͹������ǋ!�W.��VM�I�{<˲s��΂Y���~]���7�dK��)7����oH�j{5D(�
"��C�#A�הn�0�\���a
/���g`���F��)bAb�
�I�v�ڱ���DD�VG�Q��U�P҇܈�x����F�Lf(k�3S�� ����ft�oG���8�Xƣ�:[�G�rgqI�St�/�ʔ�桡�a�K3��Y�2���PJ�O�[M
"F�tm3f�(ג,�=]���Ő��j4NӔX�u���i�TA��#�5���GܚJ�$��(�^�B��\&�/�s�=n�@�a��0Hr%�uL��s����Pv��~;-{�Շۥm��{�b%֋M�o"U+��@��vP�!kï�R���.�]�
���`	�U�'t� q?r��U�>A�Y�4�o������$��z^4)��bc�Z�^�/�0��m�e���1\��㌘���9�2:T� b㼆�J�$3DBa�������r���I(��L=���0�'��)��ʰ_$}�t�r�\�D ���v�'�Ś+�w%�{=r�^�#L��B��UB��L6^�d���a��(��o��e%��{6/���V{�Pqkv�r���9mPm	�Αse��(k2�G���� �k���%��,�xb���l�NԽR_� �;�F1�೚#��q��^7����V��u�S�w���j����1�Gh���p�z��ȹ�9E�ƑY���+f��`�.3G���@hk�$����	����;ވ=����P��dc�s��/[(�X7��#&��Z���;&J��/7��)���"�,�*�d_5	l��Ǣr37�+��t��a*i�̢+v�S��^�v�3�7nSv@���6O�Y�c���G/���� ��W7���
�GF<�� fD鶼ƃ�]�E�3]u��>��@�JU �y��~��z�_����W
]t��f�nPy���6���b�}�d��g���n��y�"x6�;�6���v�k��$Π�FW�����Z�9������\��6����Y�~E-�K>�ٙ(��&�Y)�jj��3̿���6�s��熢_��A%h�s�i��vzF����v\:<tTL��|w��iFs��y�5�K3�y���DY����7X�\�n�]&	W��7��Dg[ �`�,v�g/[�M�:�����W��g�\z�=#�+�z2�&��0-�։','���y�q���V�&ݎ��!���Ρ����&�2k�� �M*�ut��C�N!��w#(�+�>�
& L<�R�h��*>��o���j�y� J��G���u�܅�У��þ:��e���>@��h�)�k�����ז�.���!."g���-h����-)�6�Qϐ�sܙ���zkˊ*l����4U�ʾ�5iw�#����̗�
�xz���3�&Y�h������rX������*(�h�l�Pf��v��R��E�K�	ڢ�&�N�*��s�`�e��!�J0<s�A�Ζ&2z/�i�<9�G'9^���J�M����jN�(}s,^PΔ��%�Χ����u+���5����S�Fpe�~�K��
;� ��)�8rD��!k�]<��btJ���6���޲ׁ���*�o!|4ݰt9);�ú�}�u�1yq��0�_�,��3��dW��ԅOd�1�Ȅ֯Q�@F���{�LR�Ի���69'D
�ޢi�y�ߟ!Btm�8L�|�N����;�sS&<{4:Z�8��E�a�B�4�J[��R��'\��0P���F�q�a��5�Ҍ-Q�oj����pG��0F��,����x���w��l0������}5���vAF:�&�z�Y$�F�[�ţ�a����@�:*�p��^KtSܗ׍�n���8l�xqs�C�fG~����o��l���/;�NᎣ�¹�	K"�~���Nj�� ��Q}�f���_�h+��W	+�x��V<���{b�rv%y��`�#�̖\F�l�)}gc���LU�z���x��ں�Ť�����-� �E\��._
��r���E��{�]�GG� 8�Ԭ�O�������Y��)x%er��ϒI�e�jU�Do��{LNM��'�<I��D���&T«�v����%��x5�Z, �e���$F*����EH~Y�i�#�m���%�,;�{J䵉�$-�}�g|K\�ʶ�@��~f"�;�V/��[��w�6V�3��bB�h�F���v����]�}�N���Ì�d�vO4.S��#��c�%+�t������mfw�����~�k!Js���y����Vq5�3m^^�AZ��VN5޼C01E��r07�A��fbA>T�/���qN�z�: �� ,�uS�����Nw��$:W��?�����T�W&-����	��جg�ʃ�3c3�f��#n�5Ze���y/���X���)tcyLl$� Y�s�#���.Nk��Wu�ߜx�v:���}e��C�^�K&syp�^N�.��/}1�Gi���:�?Ң�k�[+�ɜA�<�q���II�>U����4��Om�V�zJ	ӨX��DFwO��<-�O���3�C�i���Xj��Z(D�e@V�t2)�O�6�(�2������R�>a��l&&�\^���-"=�9W�(�U��s����₿�	D�/}F�����!u����p�)������§�B`"z�r��mF����|r�<�-���y���DƗ�S��?�����w�SZ�f��t�)�O��C��a��Esd㊑7�$��lq?�u0�Q�Bқ ו	re�/G������>�?3��cr'��hhDG_���w���o�%&{GU-D�7�]�,�fҠ�����e`P&�Js(1���,�p��!�|4���kP�w �@v��
>�,+\&�c���֏A"*I�_��95V
����
�Oj��,�i_�E��N��\ch9Qg�ho+ m�������cM#8��ztČ�W�G��TL�a��	w�:��!�3	�3tc=���p�/,����_-Ao(,_c�V��w� sh�3��:�H�r;2�n��nt<y��hᙷk�oTR@�w�� �rsl�����0FZZ�0U��Q�˭��;�v�Iܭve1��2�&��oW��(4 ��^�4P}��)b��s�6%���j= ��>���PuJ;N���$���)�q�Fs_y�J?�k��C�N��i����\lXgX�Q�l:&$�\�Qw��-��E�D��-�&��$�ƞ��
�z�$�5���d��9z'�]��k�3w�`y\ǃ�>ԡ�'
i#�+x��R@_��Y!�����Ɉ	�Z;�M˫�7���^�mm
��M�]�"��	�
�#��E��ҤfCRiN~p,���b����t@~�&�	C��7��?+�\�����9s����W.O��q�X&k �Ƶ���:E��?(�3�ށ	F
	WH��bV_����^$WPlHD13}� ��65����Kj��UW�u}q<k9[�5�P"�L@f�y��]v�g@���� *���a/O�z��CZ��r��@|��8q�K��[bR��eck���FD�T�@9���Fӻ����i3V�㻚��ÖO"y:A�����+▱�|b�SeCp�ԡ�t6��ή�O$���˗�G����V��4�����X��]��"��ZI����ח���B���`���Uh � qpȈ�x#s#���,�j�}�k3�oS��w.�>�Y�'�i��n�B��]3��p� ��_(��{tb��a8ᕚa@�P����MCf]_� ��\� I�%XQ�a^Z�� 2��eӎ(���5Q�Loo���:�`���BO��qۜ� N��U���խ�_ ��.q��u�O�9�\�4[����@Ώ���8���C�/!���oYK�
r�t-)��?�V��k��n�.�k"X�mf�A���Wΰi�vn�Fϋޫc:nz�@qF�4�,��F�d�NK���9�9VML�P���J&x�P�I�ƙA7�
�A�~zJ���"Ӟ�ښ��<�v4m^(��t�����'��ĳ�m'*O�3�y�2#���nhM۝,�Ӛ�N���/�O�V �Rp{��C�;����^�H��>��=7�D�D~D��(JYP��,���'���%�C�>����|V\:�i`��K�����bk6/B�]OpL�'�ݘ���:���j�IW���Y���;����MUP��)�cVTr����;!u�,���\9�x�R WU� ��ہA/��	��_|�×��1��S�?(�lĝA�'�F�� t�и'�<i�A� �mf�q��l?zz��^^��g3K�*��7I���\Z_��5R���4��.������\Е�cyΞ?�x֒2$l�
i�tEZ�4)m��$����x����T�\cv(�C�G�A� ����3#J��{%�ñ�����əE�.��Z��]�1�oh��H1�]79���&\|��A�^G�QV������'��W}���4������C @J�Eg���R5̈́^�?it�����`�l�V�j��ku�DRX���jr�t2ejz��Pz�?�>�=�G"���"*��t�{	gy�J�iD���sU)�[���)�n^P�C%�=~,CycW��#.�"P�/��.g ���y��q���,&l�i�c�8k`���J�Gy̦�c�b��B^�e�x6�	�F�3����R�=l��OKNS�RE�u������]*�$��SeU�	��J�#����U�u�imF@[8�5̗�kP}�$\����K��X-��Ζ���í� ��n?���pP'R��Ya��z?��CA$��� �8��o8 �:���W�m�e�?��l��٩�qc꒪Hif�B�2�A�k��QN�	G��.���L�6�8omw�d�z%��Z[���xH�jtkl��F�OT��w�4�q�.x~a���yUZ��j8b��u��WCU!)���c����*��,��)���`�ɋD�MȜ)���?�4s����J�����Le~��{:I�
	*�3Ƕ��w�5�lm�������u\QS�<y��84���܍�s�F�#j��{�d/C�4�#��*�����Ɠ�J���\�/ .>	��7:{]��dL�J_Be{��6ˆ}��"l�k��i��萩iaX�׊E#�M�N��0Y�jF��3ԛв���ƕ�7��j�����/2-���ֻ��U+�?_/���TQ�����/\����硢aل�� GX��$*�K5�ʡ8�����ʧ��hW5�w�'�+���IA,����.���;�����K3r8˖�'�h�7��T5�[/$�wv� �{�@��eB�ثڠ��ݗ�t�t(B�����Fw����K��De�]&-��z~sd�ϻi�I�Ys���/�o����i�Gs�}�B]�Q��実�m����
:�����4(�l�S�5���b�ǗF��5�Ԋ-�jxA]�р��U��N������-ߙ����E�}�CU>@���
�E�Y���pM�
4=�g3�E��	%�%��D"���L�%�{��2�OA��f��)ʫ�=-�͒��;2�j��O���m&x��HD�Ou�v�/:�i�×��l�����9�%pɁq�ֵo����@��N�Z�N(~<���B�ܖ�����p�$G�{�9rǅ��H��z^�l��bw�4%1.��i$�A�~�i�؈��&�憿E�[h��)`����P._f��[�� 8���ɫ�[��<��{�N�^��D<�'�� ��# ��S`s
c�Y	Y���@J�իQ�*o>�P��	r��7��QOGU����T�Z
�5C���|Ά7'S�Ss���]���=�����X�Gz�4�	d��"�w�[9p�y֍�G,���F��ԤU�Cl�������.������'�
	��?�Z�R@v�_�	&�&i@9��oV��nޮ{���ǁ׬!���s��l��J����a!VP:��Li�x_�9v�<�uO�.���;  ΃��S���L��4�9��!�m�(N	�_�mʳV���J�b�o��e�l�߂�����c�kW���Ԥ�"��a�
�����a�h�q�?!��V�$���,Vue�\��c`Rح�=x�,��0�Ѭ���D����o
 e?�v�����W��Xn���=T�D�J���6���")]ޚ�|}�O+�י��{��V,T~==��WB$�J�$����TQ�X�H+�B;=Wv���&���<�ǈ����>��e2Y=��YQe	͢��3F7qb���!�|�@�L�9ZQ�:�J�Z�_�tG��B���;۹��6��Rfp��������׿������vII/@�c���j@��tӨ)�R󧳍��,�q(�軬L(��\�I}�s�	�־��;]E��U�����e�]_�*S��eg�G�F�Ĵ��i�����`�m�.,�����v,�Hv�Pmb��(?ؽ�bM/s�������o�T��cT��?��?&�i8������g�K��wfwk6uؗ��m����+R��N�yy�{S��.TM�v�-{�X��E^�YG���CM�cX� 	U�=Hq�l0�c��߆�B5�L���6�(���-3d��[#�\>d�Jڵ��A�5�D��Vs�p�N�*���t�K7=Rk=����Kk㣈��4F�oQ�L+B�ǳ�U�/�ŋ ��4�|L�[K�]�͘۳�P�h��\Ug�ֲT�g�;Px�y`	>�#/}�g�itC�%/<����ZV2� ���lY��D>����0�NM6�*���޿���'-̾f�nbo��frE=���ZW�U��Q�3��̈`=�-%����I�S�J�
$�}�Z|��R�����F' k.��8�����=Ï�x��3�)�^%L^�&i";Ύ
~�f�__��! ��ǵy�-:��V�!��r;JW�̪Al3!Ҏp����pB��kZi9-4"�T�b��d,��3q����Võ��:���m+bz�g�n7��a�S���kSu�p���"�H<
�^�@
U4�K+ N=v�OH/�y%UD�G*ҞƷ@�\��n�S�%�׉f��Y n����ؖ���̅[���*!��&KЮ�� H�������ph�".��F�����*U��ο��R�q�V
.�O� g�s��[�=�^�
��EB�@�D�����\z�ݤ��cA���t7� 3E7��t��G��%k�}8Dн�Հ�Cg�T�7ؙf�@��&�x����QR��'!��K��*�7+ۚTľ�o�ߵ��PV�S����,�#��8t&脥��Y	���jv��zܻE�c7�0��_�	���$�X�[����M��[�a�e$�D��͐GI��]�e����Yp3��D���B�f�W�εKI��YdA��Qf�.:
gFs���dk\��}t�k��Q�C��o����"eb��y$k��7��kXy�V����sg?|<?��-��
�#���|�dn���[sm�ۈ	d�&���C
}�cC�$&b�5�a�=�/�L��K7��3@l�Z�)��p̛����ӏ�dqg&�����\��:g�����"F`�ki�&잿�Ӛ�Y>�.�.~��:�ۙ��N�0Jԙӵ7�f�'n�;�N���{Ҥi�+w.�]�o���:9S_��]^L�5Eh,i#���u�u�~tW'g���!��1���$ �;����hE>У}:�F1]�@Um4kg��n��7�^��h��B�4o��o���M�R��b�L��w?H�����U���X�DU�(�({تw�?��,���-{���@�M�y��V����v��G��j�B�H��C҃a����~M��I;M��4�˷;D�f_`����H~� xT��p3@NP�w�ki��7pid��<쎩��^���"|X�.Z��&_��)Q�G#i7U5�����|�'�U�F�1������p�߄����M}N��y$�C�G`��^I4&�D!�i6�N\���"8B��i�gk��VH"�
q�N0���6�����?cY'�u�>��e����[N����=�\�D����oӯ7��o\쏎vh%#bҸ��"���eQ��~�[���a:R4�52��T�͢E��&�n�C@qAu�55��/�i�/\.}=^ݔP�m�h08�S�F��ω��ȕ�w
��3-�9uk&Zݮ\��4�\қ,��Ğ`�(x���`5�_lB���?���`�ZD��Kx�����Zs�q拨�k�.�;:m���j�R�V�${��k��V�w��]N����f�W�`�ע�
�
%]�'b�.ǹD9�"����~��鞼�%�p$��P���^G� �i�P���!%*p�9�H��u�,�~�����ݢ!��ht�7?�Ӈ��Bf���-r*���?s]�T1��9���n�Ԩ��Xl#�f@��P��uCM�J�����ۤk���ɝ�s���b`э[��q�lʲ=P_E�pt3?��mN�����FƇ�.FH��j��)Ԋ��$����uA�f����~?`����U"�A����c�;KZ\1�ֈ���t�����С9*O�c`W��I��RxS�4�Z�4���N�F^�_z�~
�7�ut1��}K�M/>m��I��	���Ll�h�;�����3{�ơ����Q6�5��qJ��ʝ�9�Ae��`��8R� ��l�<�o
Xu�Fc�7�dK�Q	 ��B^�Y�GaP"�ETSv�^C`-�n�����9:��5�Ⱥ%6�<$R��s�c���3A�oͅ��Wl�=#٢#(�����\�9ŶeԂD���')\�̳��Ɵ��D�o9���6�i�� ���Z����X�j�����I#/�W[;�D~��(��A@�����X� ��/$�B�rN|���j4/ݓ�@I�٫����
Ԍ/�O�HƩU[NydB���F��F�f����y�Ncސ5^5ޭC[�Qf��p�/Bc߬�2�~(+Q\�:s5���1��oU/�(��������˸���R���3�.E��Q�ntHw�@�m$���KNh9^AzH	Y�3=֬/c�9���P،�O��Z��M���R�,a�5 ��@�P$s8D�(��j�{n<|�.l
4"�t&9�b�s��12�����V�;&���7��J�b[�x|��� ��,��3�����}2;�E��L���
���`mHi�b�7�\�5���Y�58�����C�.��g���Th���hz�?�w(�u%#uF��(�������!��w�[�.�Usʌ{Y㦱򘇎�mˀe��~��ۮ�p�D��b�K��8�;�ž^oJc����&n}�����Q�������A��+w�^2�7��/sF�(TeϬkm)k�I���-Snj�~����5��\zc9u"�/�_�{��aM-��;읬ߢ@M��q��jdY<�;�@T��}�Wu�g�0!�Z��J��
ɱ����0 -��wQ�Q�!�7�Sb�8sP�r���ku-OÉ�0��竬��e$G��xL-�q�E�V��by��0�c�ܭ�B�C�S}�]0:�+�
�#>Y��ZA������*x]��ɵ/癚x[�� ����!c_��c�v̩f�-��|��pK͓�YBl��y�h��7����mv�8�QĶ�����"ͬ��@��\_�{�����
����z����_�OE
F2�<l����Ɩ��{���J[����r�l3@�N�ҡ�xZcjl�ס(d"+)��݉
�ƌ�ˋ��5�Cl�PVi����������L�`�A�9S���^
���K\���0T@ƜJc�����h�0�3o����)'��Gekt�ޣg�8W�C�Y�)7��78X鱣�~�.7�𿉷�C{t��,i����Za)��S�]Ӌ���	U�s�jw�=C�}�,ڐt�q��/�{J�7����W4;_�lӓ�Rl�4AC}ZD��[R5��q��:C,11�v�(��b� t���ć���9��Į�o�3	܎���|�L2�kKu����\*�`]�S8���hz�%7N�3��B�h�2�J� ?��ўh���Q!.G�����.�A�/x=�i܌I���Oj���R9�S[s��)�e8u�E�ƞe/d�Ѩ��T�YǴI$�3��8$�fb���: ���4�^��Q��u�H��.�b��D�X��y��f���C8����;GU7�
E��t���B��N�nrcnX9�=�< ���럇����J�\*V���= S�	�Z���W�2�A���Qj�Y�vg��%Mp�!HD��~$�;H�Y�����96�A���\�/�]!R��JH��s;��q�ѡ�_�?�L��b����j!v�=�>��C��,iG��bخ.�]x�(�� m֩��Q����%>����L� .�x��ְ�O*��g$�S̴e�V6p�6��|��I��g[Q���`u��y{�)�&QK�B��fä���#E�t�Bh�䆲�u� ]�=���I7�Wib��ڝ(_��C� %����L���Lux굕���IQn~g���,��딳G2���PiO�v����.�t�Ub�yF9�)��c������h��%�Ja���v�!�Օ��= +�L߾�^Ha�RN�z$2����I��Fd:�|(8�/``]�f
�-Sx���>��P�����y��[�#�Ĭ�G������EH����U2��@��ڃ�7�Y�}Q�L�S� ��{��FRK���i[nj+
�P�	M劎�o(��+3�N
m��Ǣ�4��[#�ؐ��!�+�h�!����?��As*�$���9��d?��h�V�#��BL9b�ڔ��*R.��Yl�P�$5�Wn�l��'N�N�?�����Xl�;*'=�>0�����[T�=QװyE �gFk�2Z��5�Il�UB�v*p���w�  )��ɛ�b8Ɋ�q�6Ĩڇ�G����U�����p;�x��9Hܝv]?��������=4xK�	���tu.������T�t�,��L@�}���:�x^��I���0�9ֿ���ɨlzt�!����}�i�������{P�[( �XFz�y:��y�2���L'���r�z	��¥�MҸj�����%�����	g���?��H�=��e6�������0���l�P���u~Ê�����d���(��4��م��n�z���kJ&�t��𣤿RD'c���xޏU?]���Y�'v�.�	hY�I:�͝��}K4��i�ΤHWQ�EV�M��(�l��7'���6I��V��ƪ{��g)�
9���z׮�x̞G���[[%{T"������!�bX�(�PH�=}{�c v?�S�'&��@e8��" ��\�%m�'�����&�櫘��Am+���YR�E`y��@!�A���3��;,��q�_�v�byT�L��E]I^���L��DY$Cήw*��L����A*���&��ZJڹ{�5�~��/���k���s<z<jR�#,v��xa��m�D�%M-]�u�������a���_����>x[ɮir�i�p��[��'	t(�a��pnN���q�W8d?3��CLѐ�M��Nu�U��i�L�\�s�d�9C�D�V+s��Y�(�OA2ÕR�/��^�^Ri%��>Ս&��;N<�頻��5�%�]��ڗw����n��l�[�������Y&U��!�>d7g �����)Y��c[�k���J���&5��G���=Y!���q�M/�i��/���*��2P�f<��{WSQ�g]�!��Y´�5�"�K�-��go��(k�2%|EJ!�+@����YQy���̸��ʼSa�/�틫���*���z��lX�.�Nڔ�+��G��E�?N��9Qױ���Ajl{F;e%3�)�a��,�K-_5Ū�C������[�D�Jy�:=�3��5�U�=g2Y�Ȋ'b!��z�vD���s2[(�9$�����/x|?I��8�6�^j���<c��h�rhC����F���Wc���"��]�>-���ɴ�C�E�V��/y_�� ;�;��C��x��J��U�ѐ� �B�||�k�t���r�;Uh��u�Eu ����+��h���d9�K�<N�f{��u�vl�w�Å���`̼k ݛ��t�@c�,շ�c�]u��Fob�l�MԔ��`}U�d��K�ծ�����HI)��8������1 #'o�wy.�J�]����� ��Vp��">�� �����E��f8X�e���l��ip+��*��Ԩ�;s�����Q~Z�e�����U�����Їε+=��^e��D�b�G���Mf*��`lyR2.����v�=����%�͠��X��>1t����{X����$�3��ڣ�R� m�Ԣ^��MԾ
oS@F������є)\j������b����5a6�kmg,K���Ij�W�	���H�;����z�YT0ԺQN�7�/@>���x���Gӊ�g\�gv��Zb�@I?��'�͔�w�\�Y��n)��tW��c$�� ��s3I�I�wPѽ���%K^�����JG��qu=���%Ǒ����4Е��6%��dr��6�]�Q@�-lToӋ�C,X�՞9!����{6�ƧSD��*�=���2\}�/jC�Ж
!��v_߬����>�}6�uA���PY`y�Z�4X�ɷCF �E1^���Tv���~�w����P�$����gK�F7"��R�p�g�U6	+m]|_�3d�Nϳk���UTv���Ⱥ/P��p���q|S7�c���K�����p�j{g~�这F�:�p�}���礓L�]�/��
'y,޹�,g7s��� !՝��=���˵��5=��Es���+��\Y��'t�ӽt��)�i��_�B���VeV}��o�����xc}�@5e��K؈C�M�E�� �;9l+�i��&b�h>�7�	n�f����1f�0Q�QK6��c'J��k� É����W���%p֡1$<p�vOLG�{7@��i� ��f�T�|U�;�o�Ī߼i���j�8]���|��B�pD� �Ʋ�o���ND�9C�)%̈�Pl���3�pF"�w����uf �?Zt��M %7~�Ώ����<>d��s7qb���� 2��| �ԯ�$��$ӻ��]�Sx*�	)��ěC��	��U��?�1��x��$UWXh���g�b�o͘�����L"�������^N.�>�F�c((��E��G�>�R��O��Y��zUB� �Ҝ��\W���CAq`�~W�Pe�aˋr%e������ P�"�#hD�/�=�Hq%�0�k�D��:3o��N��	M�HǞY�ZF����6�k�ѭ=�ُ=�s`A�hOI�F@xv��~�N����\ ���f�ݚ�E�x{�q#���w�R��$����E�7tݿ
�RmdV��:aͣ���������#���yF(J�L���}[�Q����F��0��Iu�%�� B=���:, JmU/*;�R&/� ���L00-�'��'="�y��[�TO2r�:N�0�H�AhS0JۄUc�$�&e:6xb}o��r&�K#��ͦT�3�{tvC��ؽg��ů��T�\d���U�`�
�_�V��z��B�ڬ��1�?�Q�˩��#.�",�{U���zQ[F�xQ�xb7���O���Ȓ��aO�c/CX����o�P��,�����+ ��LP�����X�x��߻���=-V�]�t��m���Üg5i&�8K��;��0&���$�ũRW����%Rp�1v���"&�	Ǧ�?�PIW�?`��aTYF��k����-�����'���O���P�}�֩�o,"�-0�+�Pʮ)�X-�ha�w�����|B�,dWyN.ϻ"1����Em�c�fJ��^�s��r#�v��=��о
���aN]�J�&S�"����mS�|�C���O�ߞ�6C[8ma�tL�y{o	|A�R�Tڙ�=�ҎS*;���7���0,�|UG �ig��[�~\vT�@o��`{��t�Z�Ji�R3�<�^�n�b}v����	^g�)	�P�y�*Ä�F_]��%��C��nl��.l��^�rfъ�C�
1�+�G�6�k��Ɓ;�� ��2� <�`P~-�?@�u��i#Y�@�\GYz�)n^��-���R2F~����h�&���͒
���oV�sN�:��Dɮc��jB)��7`چEk�ԒLA+g@�VJvF �i�/�B�N�g��8u�*M�������w��eQ��v�AC�|1������ �bT�r���wO&$b8٭�X�.�Z8�g�;�U�pCϝ���S:v_��*��W�j�sвR����`�q�h�RPi��]��II2�^�(��\x�m�M�g�c��"�w�y\�y�7��[�5 ��8��8�X����ї.=��Q�w�K)ⷩ�m �?a��8�V,_�Q �q%KT��'�	w9�ؘP�����ư$`T�ànN�A0�I�8���w���BUӉ��b�9�����W�4�ٻ�f���nE�u�	�����a?sZ}���=:+�h��N­%��x�?�1�Q̩z��ŗ|�f��(fk�c�� ��Cs��X��z�|������J�;B��!���G���IF��W\�}5�P��5P`��w����
��c�§N�{dO8��W�۪_~� "�Fn�U�SFI���аO�����sbR	dΟ��0��{�@����
R uWnM`�D,P0��"�@�����,��Ů �s�	:�I~�PKؽP�E�	�f����xX�����=��&ԏ�
¢�v;
֛�1)۳P��S@�I"ў�<��U�5�l��q+8�u���}[.���Z�Ң�Y���1 �`�_J
���<�k��������ֶ�k�y��ݞ����b��X�4�K���A	u�(�GbΣ�R4~��Sr���yfsT��kG\L{Z6�O��~f-��N�5)�l�ZS�;�:��BE�(H���ۆp~}z����&��`�0Q)��81��vќ�˨�6�n�S|:� �����U[ �7)����¿������9O��3�4j}y��Sr��}�YT�h�$>�YT���q�N�L�H��"1]���W�EŰ�2WТt��tb�>ŏ<�֡h?JF�Ow|[��+c�:6�͓!yq�L*��Xw}!5<��.Z�N-&�R��x�ƂG:�}E����Bա�x̾�xgӷ���|W�G{���"�nWY|�\��._��ϫ��}����Ӗ�)�0m�/2��%�7K�k����1���=�nؗ�aŚ�-F�ꮀ!]�xv��S<��}�ػ�ODP��K�T*._̘XL���)=�eq�o���LO�����!�y4K�vu����:���4���Azj�Y�`��ay\7��)�p�iN|,����Y<]M����^��z�/qО�"A�.?�p�R]��Ձ���I�}�s�����G�?��<j�D*����#�1��ِ�MK+���5,�@G�;�VC� ĤY3�n�c��ލ�2p����|��T*V{��RK�La�̡�n֚��V>��"ݺ~&��{�!�b:C�
;�/���a�8 Ɲ���q#h`�Ɖ?/Dd}I�b��R̂+��1R�d�d��iA�g>'V��gw�+>&�ݔ����Gus�b-3=VG�V���م����b{�e��e���u�)��ޗt�Ƭn⠗b�ې�,(�Ƣb≕r�Κ��C�C�WB-����<��j���Ȏ3�;UzP��b,�V�ڭQv�GvAf~����!d��e�H�G��︓3A2�������$38@E�J*�x��#��I{'��x���*(�޾�t��"�������p�O��b��� �>Y.�%ֆ����l%p��FC��ϝ�Zu��ho���:x���>Ҧ��1 uµ�Y9�Q"��;TV+$%c.�D|��>�>��D h�o�ӿ���!�>��)v�{eJp�R���[c�{63N cɰ�h5��ѫ<ӡCc	{ق���9D����Z̐�g�'C#��\�2G����1����I.0��w~��^�Q4|xJ�$k�	�n����⣘��zo�Q�Qɸ�<�̀����k�}�8qK�T<�Mpz/R�i'py#���Qm��ޛI�%H|�ͻL-��HGSu� nJ��SS69�,��8�E�����=�.� 5Ew�]^
���U&�"H �é ��|����L�P��nRx8��*P{	C����U�lu�2�a��[�����#T7L�ݞ�p����T�1�&-��7C��l�l�!��ӝ�2h]B̺^�sh�:s�4Ԟ\F�gB^8`���Ha���,���I\�}O��.$BA���i(|������
B�F�b�O�}���
=#�$v!�ݰ�~�hԯ	�)_�k�1\�.� ���D�h��AaXh��/��<=�D���?,����ʞ�=����`;t�ｌu-9>�.`���9��O&�*=P��t ��������� �ЗQ+�nP����c��F&J��<�7��<d��=��&j�>���FX��a��xt�<��~\]WP%'�,7�����n�!�-Uc���6.���ejQ�_���f�6�/��&����Sh�k �n��9��`����� ���v�PA�|���e�&;�NtYx�@�F����~���[�R���]�}�(�������G!ׄ�/d2ׁq�#9�*k	����s�Q��"�Μ�[*i��X�<J� 3���r�LPюF	vu�h���J��${$�t�x�`�Z��,K��{T٬]�a^I�\�z$Lwqh"����J�Q�T��� �3a�R����DpB-u���g��H�`wl���7�	�\�R�$�x�P0E�˞b��Mo�R���2��/ U}cb��T�^�[�]Z�CF�&����B�eȾ�{�y�����9�+��.3��Zҋ�mQF�4�F�k_��oEf�@zzy�aڴ֘BO�� \k���}[Y���q
���P�fʁ�J.a]��Ƚj�䚯��r��/R�x?�rXY��ߴ��~Ky7K��_$�D��&��Jnct��J����~Qd�	-O�@A �}0��v�U���Z3�YC�7t���P����[~��
��(,��ա+��Vh�����E��"��:Ѥq��H�]�ߑ����D-���o�7��俴��j�r���+L��[�(+0i����~j���<�\e�ͪ�n�/���.�Z͜�I�<p���n({CBW�`CN&ۀ�@��U�dW5����n�z�ꉑԧn��U���I�X�g��LF~�}���F�Y�����8�^��j�+�0%��Q�q'T�lK���#X�O���Y/x����F��`.���̽ڭ~�2�#~?8|���a3u�&�	�t��y8fYuz���X.uw��-3�ً�E�ͯ`nN��D��K~	��
�j�u�MB<���Y�LgEn״K~*��7s�;ujp�tD��K�δI�a�r>o���D���Ct˝���
�)S��fo"�+:JD�X�-Y*`O��f��Y,@�bQL�,Pɓ>l
(^��r#~���-���S�5-�j�y����@ [��g���"�{4\��E�������V�˻?�C(�r��'��2qTcL� �Q$����է �x1^��l��ϊ&�9}����L������-���p�Af���
�\'��Mw�A�c�!>1 ��Dh!lV ��r��%�G1K&f�24b׮N�pM:{s������.b���@d���b���2%��+m�y���'��IxU��O�t@z�a�����$���u?4P\�&��z�����ubc&�p5�ۆlwN[���~ۛGler6���;k�rH���cRI�H����r�|N��7s~�s[��F�J�)���H,oガy")�=��gMJ��9���6����G�Y�X7)���.� �QޫEru��W�~�8�*�����IOߋ@���ǒ�^%������	���:�!8;$T>#�
��(7E+�uJt}^ ��u�~��cO�����O���&I��ٶ��pP�:�]>r�`RPo��1JC���!@V'\iXL�?|{]O�'���uWKWJf�)J#
ˬ�����=�q��)Uό&��LFk�}#�W�e�y�� ���8�����j^?[Te2��k�����g0P�1$y�A�p�4�W�b�2C8�L!7�c*R���Ȱ~���J�1���on�8���kJ�s]c	��yUCl1�lg��2coo��awp��C�������6�8�)�����3���\_�+Js��-�X�_OY,u���Ͼ֗��H�]N�ې�����"��9��<�ZX2����������A~kM��6�uбP$��^�$䷆��	RݭcQ����������5���5��nQw�\��"��f�x\j�0l>p�j}���?fH������� tM�Zuq�+��NM"����'�Z	�{^�T��G�Û��~ ��&rD��u�"���
�)׽FU\�����#�XD#:�\��{+R��	��!`�}���>�Uxjϙ]3cC�N!�{� %��L��Gs<�+���rz�ؚ_��0HU
�����?�ͪ��a�r�A&̊�>�������ɿ�/��tsNB�^]��)b��c�������UW��z�S��j�f|����r�����>�"�$��#�R>��@Oj}�^��Ψy���*�L~����-���POsS�jx�g	��芎��`���h���!�A?�.:���x5Ĝ�l/T�ĦY5"M��������������H�U]�ȑ?@�p��)W���ӼLa�P�����oĪ�����$[�q��$e�cں��ms��U9����y/G�U�`�	r��T�Ѯ�,�+�����;<�q�Nox��Õ n�f���bÅ��DQ�������#-�o1
'ÔrJ�M�9�rЏV��\�!7���ؙ���ϋɹXm(��e?�Op��^��eA��U����-�p��Sa�Ӯ���O�`�)9;?�M#w�S�tv�&�}tTK2?D�����@�AW�^jdmcv�볏�����H��u�s%�I�Y4ax����Z:�� �� �<<+���pp^@�s�����&��\��W�MFk SN��]s�?WJ,�P�v`��K�*\���U��'Ϗ�e��rU<�3���������c 1��~�E�*w��Ac�4�*����e�~�K7^�%l��0p���p'���A�����Y�)�)齍�_%��ʁ}+ � ':?e�����g�%��^/��eӵ�!�%ԉ����^&�`�#=y���M��OC��N45��&��E?7rEy�#�p�����A��R��~�T�rd�=�)�L��Y�-�d�U��/"��3q0�N�_��TO��E��M��Ӽ,��
g�� 1�&��:�L�jh���A�i�h�k����I��f������2�������,����zs�a�Ω�=�4 ^ߜu�}�p�?
��?ȋX;�iu���8����e?*1����9��Wd��
��ͫ�n�ҹ%P#�LO,r�t<���gd�� �VJ��q�&�}��Ԇ����3���Aj��u�&ߊ����~�@O�+g�M�V��b[�^c�`a���	�u�ȽM�˒��WiA��j'U�`� f'��|�?¨\�-}�e] ��x�0�%�2[=8���
�
��{xN�w�Q��:K��9[L����L;�w�9Q?\���2L��0��8�f��H��Y��-�?]�$b#
U*�\���n�J���wg{S��%��)�Q�i�B9ӱ��fGν �I��#a.��<��~o,��C��@��$��eϾMM���{/E�9T4�TJ�LP���^�S?�Q.�tV6<=ZqM����a��qW��l��2]:�wj��zH�&���&PtF5�0�m��?��#b�P����T�����9C����7�/�.���Ө���+�yeyK�O��8m-�y�3�b�deG��``O4t�)3 ��#��)@�T�2�Į�>�XN���$q�����0�b�زn����	��=����Bo[���S/���+uGK8�.hO}
ְ��<�(�iry�ӿ�&��EF3���*|S�J�|-�x�% #��Y���k
�*Dq�3�B�7�Q%��$i�}�㒟�ډ�sЌ�l�8�������G6�阄a���鸀��GOoS>@�Y:�]���C��j0d�d�S�-X�O�J���6HF��T����1:ȟ�xrq��ewܞd���rE�{����Wd.BݹX���}rܤ*to����*���	_#̭:�o�(�&!~�i��k�K�-�, Bԫf��}����g��ً����Uf]�����EZ���N��l�=����vE�|����;�st�o��dy;;%`M�a/0�\Z`k���A��`�`��>X(�N�	a�L�<�]���)>��0X8!;�2����8[tM{^��D~4�5d8�b�Ol�q�.3����͎�NiW�ʝ˵�~�#$R�B,��q�� %P(�G;�;R'�q�5��Y���I���6x|��������P�DV��1<N3�Pb��.C!��.���7�p�RM��H����82��N
��va���+rV ��,� ������N~�?[���`q��!/���K5��w��QO��9�N�.��\❗�;��K?sy#D�K%<&S��� �e��K�����P�ܑ,>�5v��M�DE~&�=e�4?���&ck�>h����Tj�ս����u��@)�
�����sv\��v�>�`FwX=�f?�<���W؂��I_f�Ȁ�ih�t���8005�y\�����=54\m��A�ѣo��T$[�(e=r��V����g�\;��P�n4GG��D��(���B����=��k!bӐ�VͧE��l��٭O��&�!z�N�����h:���4�9��WiQ���q�ǟ�hgf4�qX��t8J��3KP�Ot�&F�îӜ�^l9�G������n�`�tΩ�s���&
������աnfN�0��,�D���+ػ$(���R�-��/&� T�QzL�@DG�k���<��MS��}I�A��*��s����(�fS���H�rH�*�Ov�7u'�~osE0%[1�_"���C������s����p��)�.#aC/�-��0�-|$�c�N�&Eˡ���
	����h����ӊA�'?�DwX�f�2A	碎��LS�8�C�����X���ۢLc��J�&�kE��i̗<7jA�sX�����.��W��h���%��da��o���� M���ş�ί��#��%g�j.�b���n�����2�K��vDdM�s.m�����/��|��,o��3ْI�M���I��Lo%-�"f�d5S ��\�<�M?_g\����j�N�s��@��ՃϠ�-�]Jk �8B[//���i:�ٕ�^P�0"c�jp�_���=-����0^� x2ɕ;�ao�غU^��N���R.>�ޮD�F.�}��=�} ��bӁ¤�AoE\m��G:����<8G�]��O��b����٩�F�"�	��UNm�;���,�(����Ա�;��5�( ��8��o.��m��֑�W���KaN���o�X=	�$���%"��y���|]u\>�|B3g�SBN֬%�Ԧ�?h�������b
@�Y潵1i�6i���g���.�G��B�:gd�H� wҡ��}�n��Y`��=��<n�j�q ��L��{Y��0�h�?��ձ��c���
p]0��o��!�HSl�������tc�AH�x��Т��Z�ٴ3t�I����X�Tv6H�F�m���nT����m�aq<�L�]���eXpR�i)J��i��>Bj�c�K�Z�c��A ��`���
6&_�^^�%	מ���A]���k���=ҧ
���0�8G1���S�Q�a'��X
����wҹ�O8p�zø �p�׺*�!H1[���PL1[?���z\�]��UZ'NE�Pa{m���҂E�{���c�2(��T� �2o�G�@����~�ぎ!&C�?qX�S~�*��!6D�q���[��f�Ѹ߈�[z�U���1���9/�o�,�jF����&���GY�;ط7iF�mJ�W1tݷ����U�&u�>�H�J�G�5:��{�3E*#�y|	`Ͻ��/f�e�Fh�r8-�n:�mQ���Z	���ֲ��Ï�3#���骸ж4�&N;�{DM}�<���U!X���3�B�p����2�w��Ѳo��LGΠC��a�9���K\�2a��%�HmT(��5���Dp
�T�z����l��dz�L�U�ۗ��1A��3���"FU��D~�{��"#㝰&�_�uq�O.r\+��e2Z��'B�f�C\J[��y��͢Qr��5а�IUV�`����2B�fU�OA��Ndv�� �FYC&����J緬0�H��k�(z���=L� ��C��83=�d��z���ߙ���Vj$v�8_ʖ���}���5)�ɡ@������K��Sҏ�U�H5A�g��&gON��Ak,#�o����ҙa��A�|�g�y�Х&��u�����2H�\���w���`�K�ql�5B�@.�2���67��/�f�C#P)��7`��u%�]d۰�/���󵝹�U�p����kP@"M����U���s���
>+�y�^,}W��H���It��7��-���' Hr�bAO��z����)��F^M/<����t��^BЃh <D�ti"6����a��>!���-����*�$�/�zEf��L�~���1�a1Q����OK
��#�Hד����Zl�@���!�>ndX1������Ơ3�_y�	K^_��J����d
����N�lv�@6�ks%:��+a�S�1�ޤ�$�:X��Re`���HP�4k�e3uk.���X\�*�����g�5���uF�R�i�H�\r���\�	�گ��9_��o����a��V|�t�Ά�2�F�s/$Jx͇�k����\?o�a�1���~�w�z�b�3<{��T旽`^�EK�u�*{�s��VG��Q����v;lB�RI�_a�*�&	���$��N�ը�[�p�*�%օUc&y�1�{�o3qǰt��Db	 p����$F�v6����o��w�Qh�Cjބ�Ԁv���fu�^^z�ѧҼ��"C�uvվ���V)�B�_s�'pG��( �>*Պ�g鐐a�!�=��0W��#�)��,�^\nN�B��F��3���u��u�J�~�v�=吇�+�B���
�3�I�rA+�K����A&�,�s�;·Z^r飁����X֪���]S��AY��D�U�
1!��-qS�/���1Vl�v4{�^~O����N89��k��v%�=�����<S��,U�<��Jl�=�jz����?�VĖ�;V2�c; �ow�`\�8�Ӭ�`j]m^�,ǭ ����}�0仆C�)�՝9�#�`/�et�^�?�jg}ucc棄�B |/�وG	J�Y��U �z>��T��0���ېe$E�՚�{�����-gn���Y�ӦO���a._�����X��|M���1@�"�e�q�Gݩ���S��{�M.��GA�F�Oa��rԌ�Ĩt�ơo$��Y���s�+<ڧ�ו旄��m�
_,0�Q�[3���9�H�T�Ah�����9M��o�T1��)�� Z���Yn�n�<�ĭͧ��kEp�����q*/)���^U/\t��ђ�pGJ>q�v"�0�t�%'��0�&����N����e��Q��!đ�J;�Q�WطЬa�f�]�\1�$�c���s��Z h,W��
��eEU��%��)���JQ(uz}_��LB�<J!ɬ'�v��sQ,x�<�Zj��Â�ެ���E�0Нx���+UD���SW�����tj֗Ž��155�d��������ۧ��ቫ�P�W������n�H b�q+	��G�i9B���t*�.�(3�s��v�fQ�xs	Ѐ����\��7��vTu�F��	Q'���߅'4[�	��H�ч`���6Q�ј�0�*a�m�y}nM�Sؤ� �$_��1��㏧����қS�ℵ�$-,����
xB�:G��az��O=>n=�,O�����3)��@�Z�x� �f��Ҭe��.��eR�蕟�a��X������6*�$O�D7	)��ئ���2�K
�[h�	��4�𡩭`R���0�:��Xeȳu���B�$+{�b+;��ݥK��^//��{�o��F��_F�]�W���~]�����TG�z6�)����*x��N�(`�'��\?���ڂ��v��䖃��!�@��Q��~�mt�6�3�b'�lB��Y�S�!@r�fy$ �T�Y�&\���Ӵ���IN�ȸkO���N��]fn_���g�q�"/;h�Z*{|�Z���1X�ץ��kG2���*�C}��y�z0���H���g�j��ܝ���Ulp�~�7�hd. �4�V�I��^�4>���˞2�K��Ճe
��{��\�M�@$fو��S�l)i�c�V�Ԏ{uP��BL�a��W�C��0�����1�R�[iD����$ր�>`|̩l$���,p ��U��b�)r�����Z���w�/��$������n���P'|~S�e�i��}1�[���9�\z~���9�:�؜�D�0�~z�L�8�@NA�+')qr�Ӄz���y��/����=��ƥo

��F�iD����9s���yZBΚHnH���M4`>8b���<������Z�j@���>��ա�D�*Nzr��3	�J��ذ���%6[��Ĉ�6�K��1Ӹ�	����6vl���5��ɂ��V?��,(Ư�G%� �xX�IMZ� s`���27��Q���w�xÃr�C���#�V�F�P|6��@�L�~��j�Ĺ�۝L�jw�k�ALۋ�J���[ZK�*
x����T���r�F�HX[i����:ۃf�&t��P	Gw6/�\<3~�4~�UK�|z<�Y���Jtw���DNR8!�!�Ռy2콌���B������l��Ћ�F��L�d,�rk�q����'�!����b�8�j�		��!�Ljd�3��ߎ��pN}<������8�&z� ;���=��R!�9��J��Z��ge}�ͦc�naH��b�UI��.�z|��}*"���l��Z�������lP�/z�5Q��"��YH"�f�t|0��[͏��7R�IA�!��Qj�"͍���Х}}�l(m���kA�	�'j� 1�[RAZ?t���L
:{��7��9��+������r�Ej�a�e��_d��ȳX�jQP��I�*>{�r�OC��ĕ�I(�������ɗ��x���1�G��4et���H0ɷ���2�)��b�G{}���k�a��*-"���eP�Q�����>unE������!8��y3˺�!���{E���A�}�%�U�r�l�]9�?|����e�)�^�ο�Rā���ϑn��I�P}�Xʟ��n��V����b	�Q�S/ϐ3�����0�e&?S�{�Z�e�cA���.�Fشo�fg�1@�g|t����ĨG���ާ�߆U�M2��#� �sU
-�	mFQ#�0/����W�M��S�F�c�iM�W��?��i3���|-�tAW4G�D�vK$>#ZRO���,�u�����<m��0�Ɗ4
w�:�q5ߊ"t��%jYkVm�K>rWe�=Խz1�1������0��g��Z�y%N�d
$�:��]̐���=���**!|���)��Y/G��OhH�N�4G���8K�����ma��Q��>�5@�&�����5�w�BnE}ɋG=�8�e��%|QJgW��o~���a�Ut��J�B%����E�zL����t�c6U�^�B`��I��F�}�#t��k���=><���9�q;o����2�\�1 5]�i][]ܼ�}~]�c�EG��Β��$��"��w&�~'�@���G�P���[81�I0fS��3�#���u�6���7��4�(���`{E�j��w�$`
�8����%IRͽI���V5������5�o�ؘ�8��ɋQ%��q�O�m�# q�t�&�Z��c�~�Ϙ��T���g�6��4�|��Jb�	�y&k���	�&/�8oL����z\�ďT�D?�>R�d���f�,~̻k�&�&Y�SU�c���ť0�4�s!7X��~�����������Z,�3*����Up���`��BĤƾ1É�`�ͨ������y�m�I���a��b�3�d��U��˽¿���t��q���C��m��2?n��$ʉ�m	��sF�jis�E���_pf���7����Uԟ�I��v5��S܃y�?�>��Y;���I�	��],}�.��j�H�.�/��]��s���d���{ta��W��I�&��''�ڂ�p�$`�0����uڬv�5"t9�<�h�M*�� !��i';:�O�n�z_�P�E�~��ͪq��\w*1�b;�t��a���z5n����}��g2����=?l��9O�D?
�w@��7SХ��%>�[�ؐ ������ێ�����`�4?3J�FR��C��ϰ�f(���(��+F:�^ /<c�B�t��従������*������qrGK��\���M��{����gh)Y�+���w��r��g����~y����C;�
�m'a5��G���"wr�Z$���S�O�*] �n��-��F���m��y�[,@ � a�.G������Gw�]��,�b��o�
-s{w��y�@��$\K���[Z���2S܋߱";a_�I])9*h���Y<��bT����o�ʾ��>�V�R���+@�tG��Ni��1�.�F�g�l>��%B��ȗL�&�cL�oQ-s�~���X4G��ַo��ۃ��ou=���!�l�Itq� q�y��T��I�.5@�ߪ�}	��U�
����� �F'��`��� &,����$:V|>&���=�u��N�� n����XBX��u�ܰ�<Y��U����p�u� �ҭ�`��ڋ�r�#�e�_wxH7� E^p�3��3��8�D�O6<�UH���؝+88�!�	\9�۷�^�����ܻ#��'��{�y�j����y(3p����.��(���x4�ۮY���
_l"ֽ�m��� $Z,eiv����U!I�c)A��΋`�M*3Y
�h��y��|��{��]��0,H7-��k'�]O5L�ƭ	I���?��6����ͷЯ�
�#�"<rM���Vdq��z�g��0�@�j8�:`N�aux���N�]R�>1�qV۷�_9��X���J4�I�D���f��K1��������]��Zk͞���F�ca�e�ؼ�]ޣr�ߧ�\Dn�J�(n���8
gK��|%��Yu���g�Y����5���F�]�t*���֧˼&�?<�W�Ke*
���P�I3=���Ic".R3��$�L��i���W�>$��H�:��g�i����}��b�e-��'C���tO&�lr���wa����f�B�^! r�
Bn'����m��\vi�cؠ�8T��D�qբڂid���p�뙮V��q�C��ʌiq˺�
G�NTRa޶�t5��є)I`z7�_Ѭi���#�``�)
?�^�d!�I%�YZ�>w���/� Է^q�x<x����M.��iZJ��VbP�H��93��k���(Q�,�����޷�c9'�>�Z	h\	��_e�_�0�L���H��q�&��ؐݕ<�e�d�6q�/����*	���'[�_6JWQW�k@C�Hķ��&�5�<H1��v����ZF���u�u*Rbo���	к�NG*f��:�����gS).�z�o�,j��t�]1�_��B�zz�֨t9ndetC��rt�i���]]�L�Rquk�Ⱦ+Ǜ)Qґj��Om.P� �mM���y��'5�.s��Y~�]� @?l��I�°A������\���r�#~�|<�`�đފ���������+!��!��ͳ<�)!nKz��1������1��V]l��i�3���MeO���n��\�]�O~qv^����.�����}c��b��:��RN��^K�6c�2z��
�y`�
��3qcS�`0Ŋ�-��S�"nN��C'�Zm0ڝj`��%.=z">��Z�:=G]>Ψ�u�~�kK����Y�$�e�~�ov��3�I|�)�ق���p��m�F;9����0��߇	�IJ䷡�����WV(�(����|��4\8#ǹfɛi��Pm�-���� $^�A~rv�6��O�9��o7zW�Dm��C�� �D��fMJ�B��ib����|R�Y͎�Yv�4S ���N�����s� �Ͼ��]��M�ъ?E���<��|ӒI� ]��1G��f���9��#6I!���r�����(�6t B�i��6sh�&�ϴ��o���� R�͂���f�J�|r����~�l�Y)Ci�����]�kk��� ތ0�T&���1{o�|B_�Q� �1^:��#�ߍ�.�}�o�;��V�J�eR�6���vBN)<�8����&��uU�!ߪvhl� r�+���窂�IE�y�6un����@	��|!C����.�\#:��	��d ��c�竢i�O�V�?�I�G��{~��P�2�a��\��ϕ��'�֌U̜�ʣA�hU�˂�"Q2@���56����*{7:��u�~��()��
uV<�&��M��< w��p3V�-����Sw�e3��3�,X�
FP`�Ⴉ{';�Q��!_�����7{i��MA@)æx�`K�����n�j���F�[ZJ�%~ѭ!��Y�W4�+_q��.�(��"��Sa;D��Sst.4H73���B��'����g�7�ƽ�m
>�X���v��r�������M?�<h��� �W���̹�"���o��WAu��L��A�W�hθPIy2P���̨#��ŭ|��p/PгN֣�8o���YUN|�W����eX�AT@㌟e����R��ݱ��g�x@bf����(��4ᚿ�:�mA��X�{h�@ag��g�SB }��`�F
�����c� ��c'���՜Rvn�O(�<����x�3�¯�$C��Y���7D9th�ar{�*�h�uc���!�m1�hxǟ�Lt� ~H�M����*A�^Y�>�6�|x{H"���e��ض�
{Kc?�4��)�<�.��ߍ=>ͼs������yk��p���n"|��dI|:���#u��D�6��y��O��0
94��3�����D����{Ҕ�̛`�%�@!��Z:|nd�aYq��H�$�`�k9ۗ�L��ϻ}�/)�I�w��ޠ��k6m���in�h�ɝ���5���~�m���0}ug�F���ٍ�}\��L)���F�У�T�k2�6��i~e^�����Ǭ'�{�s�q8��� h�FQ�?vQ��M���A�(������UY��wnfg5�k�G��漬+���w��̆�D�o�q�B?ӝ�{������������EPDE�J2�0ǅ�@0h�uq��x��*��T�_�֜�Ix���R�**it�ͤF,�W��r�����/��}��� ���cM�~��WtQ�;:�<��6��i[-(ϵ��>\Γ;�ro�$�{�ۛ�������>��J�7�sΞ�������Qj6�����Y�S;G�3�OLCS�S#�`b8�:]1��`YsCƻ��B���(���:@e�V���C@��L�a�l�8|sW����R�ȇy��gn�l/�����}o|��(S�}��3ͼ�!�j�"�6Z���~��­m!ވ:�}.�F��GI��m|��0+v�-S��,z�Vk}�0��LB�-4���X��a�.U����@�\
zTj&׈"ӑ`�4��$>�KH:���6)SC�ii�Ǚ�SU��iM@B��OO>Qڸ�Y	>1+����0E��i�����0�VÓ�`A�"Zj�ݮ�@ٻz]H��`���?9�h�5@☨���1� ��!��$����Y��I�,Ui���u�O����`�ҝ�*�hqo�
b�5��Z�Q�-��DQ FM2�Q�c�A��	~4�F��_x�_ޏ��z�(~L�*=�@	��e�Q}a0�5[/�Ny!�+�"dS�甄�0�!!ԷKM����N8�gF޺����OSz 4�����og��3��a�r�-�A�W�������g��?�3���sW,^�eQ���	ꎰZ�
]��<�YY�'Ǝ{��rX��4fpD�����!}u��(�����o~�]�Xk�s0ѿ̲_�'.#�m�#���Q�}�p��SN��s"��ݨ�+6�B=\�
9��*Λ�X�ˈ>�]&{|?��RP:�|BBV1�=�mBi��om����Q ��م�b���/۸|��M�ߕ\��[�3��Hy���q�ӓ�$�������vV�vo���sn��}&�5��0��4������l������j��<vC|�p_u ��<{0S{���p��Kv̨���PyP�6�TP���ƕD�} X� ���`��y���q
m����vW��=�Qx@��(|� i��qp  �h�Ƣ��j'Q�r�Em��n�"	���z�tM�hxjV� �M'�ҳ�fZ�
g�_7lT��)�_{�L(��_˦F(�C��:R�$�W��%�jFq�e�q���������M�F���V�rXZ�z�T�L��Q���.���n�"��6�ly��Y��M� \�Y�ū�]ٮ�M�2��!���|�,��L�<Dk�/��[l��@%�kmΐ���e�NU,C^���Qb��ȯCJU��h~�km.����W����'de����#4���V�,@)j� �7f�$lv�!���&��T�bO��Z�Y���&/\o��L0��8�gO�d7�u_m�{(����(4�Wo���Bm8���&��H�7�����'c��u�uɊ���T���
�ӟ(�V{v�W"��oZ\UK�� �\a4�F��4�p���T�`Կ����R�!�J�5u̳�<м*� �w�~���y�¹��#Q�m&����Kt PO�{�Ĝ�f�'��c��>�.Z=��|vB�s���w�A�� T�mώ����ҏ����	���yA�B�Ԋ�&��+"Sikہ�
������B5z�h1p�B�g$.-r�u��5�zm�p+ʵ39᥿F<�	�z�r�P	�B�ҝT>��X�N��.��M�a�;��hVir�Rm���y]���d2ǉM,�~ة�4��[AI�����@�'~��N���
�^ϫ��h��J|�l'�C޼U~�|	�~o�3�sZ�Kf�dY�z�Rw�����������jP��8�V�I���@��6f�g��L�V����$*}j�ɿ�<ebߕ$<��M�G㽜  	)54�ՁB�m�:�C�����t]���Pm�����&¯"iM�r��Oc��6���H�����}�vҢP�ݜ[u9k���6(��>�hGF��B�[�S�Hq	�b����>ݥ�E�ϸm��x�w�w����$=ԅ�x��k�$΋�l���I~с�� �FYV���*������@�W���@�T?��>f�g/�}�LՁzhw9j�����.4��R
�2�Q�aF�J����'3�=y�9�1͵�W'�D�31��-+3}�C����k͸���^��Ұe�tˑ����3�,����|8R�dI��1�ti�q��C>P��:V����ai!�c��ԖG��"�v�)�� ��6w7),XG:b�yWk@CX��jx2�<(�F�n���g O-H�9yZ�g��ÏUOl �ȄW��}��c��_�	M��{ȅ)� ,k�Wr�=�m��qet���U![��t��Y��a�0�Ս22���+(.�ntRZ;7v�TA#fX܌{�ńE��Indv�2�w:-�J����[�PƘ{�)f@%�Yj:1����ad�fF>�};�N�f��]]t $�z�����;�d�|/e�2���:�$e���'�=/m�R(����D���u�XdO�cA�Ws������2��8gY�ˈ,�dNy_����u��1�r�R^!F�@�W|�q;}�yp:�Q���c��(\�����Y>ki�b�?E0��������J��po��Q*^�E�0�S�)5D���d`���8��?��#'tiC�+�/9�/�+��}��>�H(Im�|X�[H�ȸ�F7/t�1O�K���s`����V���\E,�>"�%�N��n����^�:�*����g�	n�tY�[�?��I��T䄙Δ���"�#��Ʃ%ޖ½Xc������Xza	9n}�nDZ�w��6�ۦ��oe�@�	���Id�=!��l���vm��W#�w��rH�: a��� GK��Ԍ���\U���L�ǡH��$Bf�7��U�V�S�=V�09���7�H���O�ˎY�UR"VR�����ew|�	�X����[�/�h�d`�j�Q��U�]d߶�n2��[���� ۣ���nc�P����o���S�y:��:��En;��+@ML�M��ζb
���q��82�*�[���T���8�L��<��ДE�K���H9���t�Y
�k���d��5����]"�O�o}gk��ր�9��3	�?������f�}��%��eD*тӔE�<�8da�$�/̬Hu��˂����?nH߱��'v	7/��ԞE���R��,rJr�/���z�ۗ�"̘t���Y��V���YXJ�����F�=�W-O�v��n���.a����Y]Vú���B%�o�3+��M7,i�o}�6Ⳑ۩�IѪ�|��s@*G��6����v�\&I��c��A�V%)���xb<��LA�%�U���R�?��cZ����ʄ���R"��G��ʂz'�4O'"* ��EɺS�p���v��o����"�5@K~A�T�n����������Ej���;�pأ�y���@�:��m3[�W�j�3��t��1�U�����a*Ho��T�n�D�"����X���j�&�5�9u11U����;pW��kU�/�p��s�`#���tC���D3��9�}�>A���x�ᣭFm]t"iWd��1��#�>����� |�nv�z_�б�!�U�xe� /��n�9�%8�O18�=�`G���s엻y�L{��;�����)��WB1t'��)�c�ۡ ��[D=Ruf���n�DR���5�<����D���9�:gd7&-�=��qB�I����?],ێ�~~���.���c�jsE�|�l�e��YJ���H��m��ɇ=�!5�L��G��!�����0;n�߇f�@n}�~��>�g���:���y�7�l+I	�Z��D��y�XF0����N����e��.+T�N�L�q*ٹ�����;�C� )l涹W���pGX	�L�����֬�:�H�{��l�t�y`�Tj*^���3/t�	`���P�����@!�����1_���E�P�WS�7 �(3�B%Px��q(�(�c~:�U�Xc#IL��~\��2+��9��Uu�mN��
������p#�٫�r������%��:�?�+�MN=8L�.ҰXLcS2q�[�h�YM�ڜ��2��b̛N�r�c�-��:xo+U��O.��h8�����B�~�"��^[	/�gu�9�I�l 4g2W��>�S,����e��{V�1��[~x����}�����np�}�Ɇ/3C�OJ������ƍ6�vO�Q���;}T|�y�K�-��n�$�Jh7��L�j�O#�mm{9?�)_
a�q@=Q}�FETyW\^+���m��Kbv��va�b[��ފ���C���9�*�����ͤ~��e�c���1����sqg��{�i�@��K�$)�����R�_N���{���x�4XL��`Ѵ[F�+Ї�ח�����"_��+.=� �R�f��	�zi:�U��I����������
~u������H����`3d�����
�����4(���>� ��]|�n���0:GteSA����l�1������n$�@�v5�v�9w#�%����z����&�ǲ�\a��(WYIu)��gA ɞ����X��4[�������O�4"*���K�����(J�J��u�&��P �Vv�׊����XF~��-ȴ�삆���j+3C+�K�s�L��v	A�Һ���-���2��%먝��
J�Be��#6m��Ӽ��v�%�jG~����n�2�[��i)K���-ϳڵ���P Ŧ�6���g+�P�G�Eqd3h���d��6�\�'ª�D�ʜ�(�p��3� n��}"���@� -�)����F�~͌���LesdRF�(�]�̉Q��?��ĥ��OȠ����H�B��K��=����ݲƄkqo.Za3���x\����*��% �\V���m%��cn���I�m{A�|]��˿I�x׍n)��n��Y(wҀ�;zNe�~8�)��D�P�9*M�]v�Z���lEP�`F; ���f�4�ܜ�Z��h�)E1�{��i��O��`�u�j-H���6B�3�ǾT�d��+b�e���'�2�x[
�:��`��uυ<T7����7�|�1�<ͥ�5Щ�r�w{*�O�ɱ%�����Yxo=)Ǖ$�qDP��<��-��rbe�r�Q�,T���(���~���y�#�Fb��Z��i5Y���YZ���@ �U	7f`�6_�gh%��ǰ�Gcw���.���QA�et
�G�b�GC�f6����-9�4����0��D"�&�U�]jX���e6�(���DP�l�+�a��r.0��:_�9(핼�!�����	�j;���N��=�����?\�{%}��wl�%M���|q�g+�j=I��[�"��Uz^Z�ٻA(>���`'����B��jH���k���Ak�ɝ�=�)5�1�<O�S��c��;D�������i�0�˱�j.��ɚa�Ɗ3��,���{�K��-�9�SA���0Un�Z_R����=��;�I����tg�S�&���Sf�)5�������{���$_}zd�؄��"�쓎+�-��%�eKG���ā׺�T�1�����Q_p��I|��Ew|������a�.�i���cq>*Q�|/��}�H��i]3���E�L��.>����
m8���0S��W�s��*�Q��B�� E]�i��O��"���"��p��|�Sc���i�R��h��}��ލ��_h��M���S��wd�m�X��l�������e|�YIZ5�a*�������n�� �C��.A���:>8:�3!J����r9e��9;I~���Y��q�i��خp|93z6Ҝ��y�\�ў���ڬ��:��q= ���cq�̏�]�Joj��N?/����T�Gm�(T�&�d�р�؂G Ȯ�����Z�*5�G��S�헆쏗΍����+�X\�7#��GJD�
��)��VZA2f;2&��#]l]w۱:�8��o��YSR/�Zth�R�9�����r^�F��c��	���Q��Ƙ ����f�3ʆ��ǮE��@��M��yU��զ�Au�����>.w+��l=�M��M!�X�
F���BY	���h��@�_��~Y�]���y-Lū����P��Bv��!�#�Y����츆C(� �00��[ew��5�07[��8�-�ٹ=+��.�(���P��'{��|%֮�([��D�vĄ�	���M���Ƅߜ��e0b��v�i��㨋G�R"�E�;;o��f��l��$ÂjmZ�/����o�`�6Z�E��
�p^���6���n�ճ�sb%y��c{�A���;��
Cp�r(�׼�V#����N2hv�ʜ k���WC���Jך����ޠֵ�^�`A�*>�4v�^T8T'-�&�s�d��1"=�u;�(��Lد���T��#����ѓߧV���h��������h򠭿����MǤ�Ɂ��	���,�.jC~ҀkR��?��ʫ�
f�<�]��0�6C����oI�$��S�y�jPk�[ZCo�F+NW�@��4դ����;�^X�[�B7�L!���YԖ�y�FB�[_����=n5���V�-���<�K�ړ��m_�+ '۝�A���΋�6�}�������oKi���=,�̽"W��*��{��߀�q-���<Z_��b���=kqjzŤĹ���̣d@��:^��Ł�I:K������'��h�ޣm;B䰳�~�<�ۣ��A_@�	>��"�"!���;7ZL~�����������]?�=������ν�A��ӿ���r��L�0<�,�Ɗpb�ow<+.�ֵ���Jg;��}Ө�f��ɛ��[�c�_/��&e%p���MmB���M��;x��\/��jk:/B�_jhr�Q��)^��iz��� .�]�_p8_��&���E�LM %A��!*}2�0��O�eT�7���ȴo��֚ځ���k<�.'�6>[�|�x �U8V.f���J�-�@Z#��h����jIkut7��o����&���xL�����I����m���SLJ9h�*��
�vy^VLы�]d��~�L��������S-�@����Bz	�G�,}v#�i���Zd�|o��*U��Y�<���O��,��X�h'�;�O�RP�ˌ�q�	-ă�V�"�V(/׸��W@d�j;���$�Yg鉀@����Ϸ�\���_V�]�󙨲e	{"���i��;�\�NƵ���o	%:�9�@?E��p� k��YqZ�G<�81&�Bi�r�c~��=�d�#�rp'Q3������i��`E��p����(My�7[o��4��D��g]�@ca�T	��&~��I�ʖ`}c3��Z#T]��q���Ap��q(�;���a�m�YK�4I�I���7 V�ѳ>�+(�!���|�m�ZfZ�č�U�����|-�l��;$��u��$�ȁ|�a��@��	T����=�2��wȱNeM���18`D��n]�Nls�C��l�/�ǜ�7��&\����R&�/DB�F���e5B����9WM�Eː�R��7���a٭p�n?��~da<��6wn��r�_�~��Y�X���e��(*Y4��.�Z�XYl��˥�6;�x�,��/'��U�5���DGF}��a��X�q�P�\N6��p?��W6��p��K6�vqfo�6�vG/f�Z�� �8��y4)X��Û�XLͣ��!9��&��/Y����b5f!�w�����n�=�����a}��Ggp�[R-�Z�MU��w�v��
idPW�h�E0I=ï���y^܎{p�Й�:-.���� ݟ��X_�Հ)8���L�(�lű�D���2[��w��0Wv�|��H��դ�Bi���I�=8[�-KgL��~����R9$ij2�������i���U�X?a4�*uS#��,Nl38XvGI2�7Hg��5b�s�n���H�i�D��ݒ�|��4���~S�8�,�.�3����'/�՟�s]J��, d(���G�R	I��(N�*�x�`�G���)�o&i:���t���b[�!*5�xh�h��ǧՓp��nwb7������hU]���-	������&�d*����ĤZ��W�}��-:F��� �@�J��^��^OAǵ�5�� �V���A7� �|���M�ȥ臓)��bq����E#)�6���e>�y��$���t��l�	O_�����z�h_��C�~�y?$���]�a���j 8��àA�Nc/Ȇ���s�9[�sl�)�o�Q�����/����®Md?��$	� }k�!&AwQ�<�4�2i,8YI���ʫ�HB��57���v���0b����l���*)fdJG� gO�IG�/�}��MwI	�OX� �m��s)��7:<3GWR�!e|g:���9{ up��E�x�\Wё+��X��%	Zn��+��������YD�x��7��g�E2��Xh}a��2�MLGکO����:5#L��tOs���^�`+���5m��3��*w3ʵ��I��9���.L�aiS:m�E�}�= ��K���f��#�@�^X�e�O�afoz���<��Ԙ�'@��ZeҨ��8��M��y�~���f���	���LJi����^R*E����dR�?�x�D/��%��Y���n�/n���߁Ǌ�'q��,ɷ*D��MF���Z�n���e#�x�W�w�Tqr9�̄�B��8!ը� H;���
�4�1&Cw�� [7���P���_��IՐ�'C��f�6+��je��=�H�?oӵ���6�[�H5F�����m�J�5�O��A����E
��i>'ImWMp����,uw(��r��=�)�yt��K9���/f�O�A����=ۉ���J��L����4��S7�:E%��xwЎi��Mk)2�ν�"F�"�����?���כ�^j �ڄ�y "/R�0z��[������ޥ� Wz���P�7��!�F�Mn����aP!�ˈB��*�հ�D��K�:GJb��)�j��/�>T�y�?#�V� C"�7u|iU�#���R�I�r�����eZ�Ǟ����L�)A�@�#
}�����s��w',���O�*�=������q���<�lsi�������g$/s8��l��l@u��u�R7�D�+dO�M���ሑ����`���n���C��K��C����r��<u�-��\���p��M� �y���Gп^�XE��8��\&yݩg�W�/����Z�x�:��D��W��We+�ߛ���=I������E��������<LR������4�l��a�-� �_>f����w�E��O-^
Zu	�)��z�,LY/Ƈ���[&���a�75�bMm����?#�ʻ�l����{p?��={�t����'�x(S�;&�T�8nlu������a��[]���i�^e�Q�z�����^Y�U|O^�ȻN�N��|=�qD|sVf�*:!Z�Oe�۬8f:��6��vT���+�/cL0
�o�K�sHk��3�ʬJ'��Vt�[�� �#@�]��TĜ֠ ��+G��w9l
��Jۊn��l
R.�\V��8?�ߟ��k)��ev}�ds-�ن�"n��5��w���K�/��Sߞڹ�����=�u�E�Qe0v�ZK$���ϲ;#�
��e,@�{0B�}��V����ϥ����>J�L�>�Ko��c�Ð���IB��F��(�)�mv-5��;*�e�fA^qJ[!��j�a7��J��v�����,�/k@�3M�W I�ra���/
�'l��,>�g�!�w��R��f�������.�;d_Y�af�\����w�Ͽ(8�S]�����L�P䋌��@xeRp=[�a�ፋJ3%)��î���RQ-M�9u�����C���g�>^�5�Ի�'��r�/+R~��F�ف]�Y�w�Y~�t%ܤ3�;P�>�`��-:���-W�A�6 ��l�/�5�)ıv�e$�/�Z>�*��Z��I��%N�%�K��rF7�,^�_!�S�:O kĀ���<�`
�GRN���W��E�ş%剽bا)��@�����Ɓ�L,��ʼ[�&��W����B��������.Tȳ��!�[�o�k��?���͈�E��Z����GC�t��)�~�z�lvqn~�%]`��X������v� �m�/ٰd��//�����Ο�Z�c/.�j��3����GgL7G�5��8������H"E
�ե��kU��瓒�w����y~Y������v�����pw咪O+�P�S���Qܭ�7X�>y(|��n֐`���-+�8!&v�07�A^�����o5̻���S���J|*~�G]T��p~���E�
`Xne��h�u5q'��`X�<EI�xU�pˇZ��Z���7���[��������߇_C��kM��@i������T�M��9��Om3A�+�uJU��T�����m_j�=����: �1���۟���c�/�&���iE�~��kz��>��IfN1E�#Vh�|*�k	e�>C!�%����e?[�Q��B�Ƹ�޴�)D������zE�Z���MA�`�4h5��-2$�s6�צZ�dCé� 0�d����t�$�
�䙉�X���X��R0l���%�0K"ЛұM��=����IE��j��_�ڥ�6c���|��r��vy�r$bz1�ˣ��N-�L�iov��<z�ئ%���ǷLL5</u� ���UDXť�H\��!�t4�0~=��8A/�;E��Q��/Z/Kj�Tz�"J��C��K�sԩ��{�#�/��G�a��V�}��3�A ���x���rdgfO`����l���㏇�h���$g_�h��p���R��7����T�C`�(���;�B�����x���k�,��%$>^
�/�]*,�84B��T��߳��MT�g~���bA	ʼ=�F�����;ۏF]�E��G���/-�&��s8ۇ�N���Oq+Vd'�>Y�@��Ώ}g;`K���ql���	+�܄G��$��J=�}Q[�����~l���I䠂ֽ*%��,t�0�0 ^/j�G��]q��"��P�1�EoSn08O��.�tӺ;۾h��+f�ʌ��I�o���%�^�b�[vTx��x�H��ܙn�ʚʯ:̢߀]�.:',�r�
��Q���XB#�*��L.x��W��T+���m?�U(0���?���!nD\|__�x%隊'ҶW�JB>|�\9~d���s��Q-���ŕދ��ͳ@�k?�^�o�@:���S�z��O�
�Yʒ�Y�XE�ήHP�l�T��0�Q�q���
��� @ Mꦼx�}�ɽ��(Qu)���������hb�z����=<@/ �nT�0�,��֫���v:�ޑ��K#��:.�\�`��?���)⮓�=����m7��G"3(��S��n�S�=d�vY����As�-s6>mR|�_ �IS���y�������ch��Mm&[å ���cX�8�[�v)�Ĕ/�e�|�+0�V,�Z`�OӚ��<�eJ��$�2��L<��a˥ς}&�(��R�3]8J%9쇝�\`��Bo����V\��
Q+,+����U��| a��_	j0��Az�p
*7�V�P�
;�z.ux����l �އ؎	�
מ�������E)u<�F��Pi�%��Ŝ��U��<Y�l���$��m۫<�s��=��k��'�i�e����e~Y����^��Ze�z�l�_��͠!�N�(�a5�y�j	��
�fhf�5=Z|��ks���("��� \ʡ���X�U��^t�oƱ넼ɨX-����Rqc5����vm`�i>�j� =:��y�$��y�	�R����^!?�'�?�YS$.�n!������()s>O	F���NaR��BFy�ng�EZS
�_c��pt�,-�͇�f�^<�<j竃�[h[,M`,�~���W���?r>���Un�U0b�˔�fsy�b���Ԙ�T��C�G�����y*xv�R�U�)��6���ZD�ǛK1
.�+������w�sa5{w��3(R@��B��[e��ф�0TP"��gc�90��T�k}��0]���gi���$r���x�#�= /�<�IB�_������{C�X^��5�$Q~����ˍ�(j:%�%��[�UKX�f�,c�9T�I�[����>�v�a���`�^�93�`�j��v�&��v}��p;���#ɡ�4 �*Yщp�
�9�}7��B�_S�����T�'�BaXM��~k0�CM\}s(w;}���`�����������1�"�(� .2>�e��0.�'~�MG��W�9�yu�2��S���1�'�f(����<"y��t!~0PI�l=�m9J�~�z����O��"�+ct���1�o��x!T@LZ�
 L�ԑN)ի5K�A�?WO�� �:%)P3>��)�Wl���qM�PTv��N���ů7@�_Bi���t���Ռ�Β*U����x+���u,���>֗��.���������}���J�
;����H��gx����7l@���BV�s�lU&� ����������ρ4��8���N2�"�{��1T���!�Cb`jEe�sjĭ4��w�{{������<�$Y�A�^%��@�z�D)�	`�"S�K�GЊs�O����� �]}��d:`��\���]{kR �
*�ޮ�� ��v�Ty�#6�ݔg���E[��50h��H0{�|���7�kX*�2�S�K��F�-���ޚf��J�Eorb�1[�����؇�7��ty���p8.AS9�=�\�m�P�[�����I^ eC���V{�Si��=�����㊄b��.8�c�RP�q%��؏z���n闠c�#��a�N�����GԚ��ADc���G��Q�1�s��h�Wq6�%&��~�fv,�W}���a�OJ6$�>"#4_je���v�P?���z��$E�}j2���Q��U�e��YJ/�_L�Z:�o���p� UHa#�ߍ��K�M��߾�y�I7���{@�?G��}��9�	���{�[\�}� �t̿��?���֡�>�J��n#�Q��F�gsi��T�d���S��W�g3`;�-��Iu۝e�<d����+�`D?[�*�}�4'ŅC����G�a�U�Md]gu�-�G�u�xK��t/�N�ߖ9���"���\YTm��%�5<�CzC�<��^15C8�/��Vx� ��f���:���v�<x�f��k��4U1W�Ϻ����O�zN$u�e^W9���L�<m��!F�3u#^�t�;��M-:R6/�d�%�
�0��jH"$cۿ�Y;�t �����ۜCh��3_��s�Em�S��µ�ou�yS����z�x�Qq��dr\��F@�IO(�B37��XF$�ܫ?AU¡�=Џ��V��,Ɗ;��.
�Y��E�9Iv���\L[���ڸ=�����?���M%$�H��f*��+͠{�".h�*���$�{�D�6�I��/F��c�¤���
�T�i(`D�D�<�շn?"V�)|�%����ip���ڏ�f��xc-ƛe�6�ջ�����Z���s��| K���M˒#"��YP�
 k��a�(��%���MD^��Z� ~N�UR�n�҆XN�2o�?w8�zo��O`����{�����n7��FGU�j���t��1�54���L���|[�g��ZS��}X6��:��z"-��\�:�}W����dX��R��Yb�z]�c?o�a�bsK��}���r�����Ъ��*Ybԗ6̘�Dy�������J]@[���3���w�~ؚ��;���OL5�R�0�5U��	���gB/�@M�d����.pY�'��x~.t���^,����Kz��P@ӵ��]l]㋷��&��\ ��e<��А��Q{� ����'g��$P����՝^���=V�^��o'\U3#(닟y��fV��)��O��A�O�M=��/�V��R�S��~�bSb������C�	�]0D���Ą2L�	�������7l��~��K�����U���QG�~�^L>��$"��fRo$&wˆ��wM�G}�F$l6�g"b���P�Vӟ���L
٥�î�����b8h��^���i����խsu�m�!���6��D��h6=;���� ���4�xF�C�y��	�;`��!��a��{�	����ij������y^�v�|M�� ���8?��GF��v������)�r���:8�lv������N]����Ɩ��n����B*�-\l����g�>�]�P�)?�_n�c�v�V]�i�����A�I��H$��h�YdEɄ�dlp�Cpp�����@��Fl#}U��cY--<+���Nt�ʮ�5��
��N|�	X�����X<�^�#g���n$��ZP��>[��Jb솩#�ЛRڇLF}G���klg	Ǽ�e���t�Ď�}����G��`%�u�$Q���U0�\����+�G.ӵ�Fr���$�7��Қz��@l�>.V�Z0��:��?z��@��([(=�T����{%��Į'�Mܽk�\�hNy��F�Y���� ;�;g�,s�C�TU�:@n�j�\ZG�����SaB�\�Rn�*I��J��ՐY��:v���x@��O<����y]ګ��]ص�p����	>ڃ���
	�C[ ?�$p��
nX#X�1�ͩ6��;�-�y�� :��|����9w�~��}	Տ��|bu�+�,�۟?�5�0�Ѥ���k��:(�/ �1�W��f/�?t��rxZ�(��kyKG�F���dW�۶�S�-��؂��.`\�ʱd~L��f��\�kT� ]{��wOЪ9.�0�F~��x?��(�3ag.�	=�g�a�g��bfr��]r�ˌ壤�2w$���ݒ��W�lz�nV(Ȼ�(�~�3���M c?VJѨ�!s��V�	WH W&fz��;L܌j�-@ѓxc	
���Rr�y��~j
a<(w])�!��A��� �a����>�Q�u�����Z���xu�?�;? �:Ūƕ6��;��$-�Z5D���ɘ?����t%��<�P+$���2|2�d+PGG5�s>Î=��'�g��s��I�IYr��J9R��A��1^���}�B|*Ȱu���8�^@�	�ڽX
�olRc_^���1RJ;(���IWyDw������r��N8Ҧ��kd_pc�#U�M�?�����64U�D�%Q!$F`� '�b�~�aͬ�9�XH�-��ե=�3�:{�!Nχ��a��fs�H�����	�q�\��UM���?���p��{�a���Q��{¢���.Fz�����=:����z���AK"^VWQB7��]�qoR�(p}�c�uVK�$���*3v���VR}�w�~+��:,L�>��8T����v�%W&�R��|�u<e!����Y)~��E���P~\���a5�I}#Z-����>�@w�����?�����WC�힯v���2�-�����2�<��ǘT����v��`�~3t+_�}KkP�3<H'U�����a�s~*�-�9�Ț ��������0FI���V��Nw+�K�s���\H7��r�gB�;��x�?��1�XJ/t=�V��U��틺�/�S���ӝ.L�GR��$�N|$�
�o�R+	�B�:�F�V3+�ڶ䩇�x������$��&x��]�%<��ɐ�X���Js�u�ic}$�C~����dOE�� �ʰ'�}���9��^���ڼ��JM���䭋�r)���-7<m��×�K��N�������³*�H@ѹ|��G����uxm	�T�����'����+}�������i���W���$�>�]o��*��P��o?�</���<r4$7:�V�����<n���z�c�Oc�በ?��j����!����P e�c�4�e�1~�օҼl�`S@M�,�nW(�'��T��h�$��b�Q������Q5���^B����~�;�g���Ｅy&Y �� \q�ɘ@�:s]H@�sl1܉a�Ok����-��@�mF}��B_pb���V�#h,��LԌ����J �����^xٴA&��
��\�#"[{�b�v���
>�ۢ�R\�w���ￖ�Zǽ˒��Z���5inr,'�R�j� �ٌ��-$��9�e��/i!����x?;�/b2�L�fإ)�0G�+
�c��V�505�aF�|�����������r4s�ؙ%s��?�Ϻz�p�nSV1���X�Ʊį᥽��P*��}��
%;П�eH�L���k`W��SF~+��bL����m��	�-	�D�p��&1("4�ӽy̠d��ڤ-9��|��O�#�j�A��fA�t%�et}�&ɩ��]���hx\#K�Q^O������(^SO�EQR1?2�A	6@�[Q"I��3����GR�?�oԓh�4LnI���
#Ю�7S�y����E���+��z�)X(O�����)hl�vD��\N�Y����ۇ��_#��Ufˑ� 
ke4�A��n ��D���Af����D^��_20��?��,C���e��޴�(t�G��|�1�G����2(����Y�}����ܒ�uO�?��M�=��������c��-�;ي�JjH�J��.S(
Cpx��d�&W=�=�"����)���3w�,��?k��g����i��fܥ�;�z��`�O��XC]���f�7�ҙJ��e�aw��1/-.�Z��s����CH��A�!�,ɐ�����W�󻯕Mye��Ѩj�R ����f#D	�MP=����䷳z@�m�C��LO�v}>pz��	�VU\v��-������X����׼;A�&�1, �A�p�HI;�Kދ��`��+�:�	���;V)�TޫĮ���N�����S��9����	CT�(f�g����i5��N1�{�����Z'����	#g�M�8����l��
�/L���5PЮ*4MK���a�����d�����T�qܲ<����T��W�����~�sC��B��ݯh4�E#/Y���(���*m������~ܝ>�H�4&C��u�Ƭ���T�A�^Lg(�EE������e7� ��MPn�)��&;�}��:��7\!�|e�jd�c��)5� j���/ {�Ax��Aƽ����B]uU�UРJ���j�2X���&�vEn���xt֊*��|`'"[�M���G�=�����
&E���Ѐ8~DY.ÎR����c�T���S�c�q�g�D�X#���K?K�
f6xa�����`9���$�kc�4Z��?L��r]a�I��򕺆̑�<�Nx�XT�b�Q|��n�Մ��8jT����rq_�|rn=#�X�ol����FG��mu(l��6�� 6O' �6��x���x�QT0n�Ǐ͵|'�{��G��}��F_�\C?5�_�1���+h܌�%'�Й)HP��h����Z��A(+��(8�L�d�Z\���k������Bﾾ��&I['*;��y�Z�3���̝�bo���T��Tl�C�9/u
����ވ*W{� �:�Ѭf`j�y�$����p��Қ��g�����̰0�	[�%�{gEw����U>���q����]�՛P��b'D� �ހ��7w01�y��Æz�4�-�w�D����V`#�߷�IꔱtN��ܶx�H�cH�3Ƚ��vUr��K#�������߆���&�	s�!>�xH� ��ΐ��͂l�P#�<��8�*�/ty�Y4J�ɏ�p�+�YE'���?#P���2��&C������c��0����$�^��Y]VW�Ļ�\��}�˰n��gf������0?�j)��bo���	pl��mlH��/j��D3�F�F��f	I.%hT[��w�NϾ�m3{�KK���ܛ��~S07�Tq�#��e%�F�����\t@���[d�]r��_C�k�Ǌ���&�Ʌ=$�{�)���u�b,{^rG��j�B}Ukz%rKJח�rf��T�R��>*!�v�/�˵��W�{)��(τ�Ē�-�w�H�ӴP�,��C�\J8�,'~��aAŮKE��jz���|.�l�1�`D--'Hk��C}��"Ǚwq6�
_��f]l�L�^j�ᡥEk5a楤#�Q."tq ^S��(}���,�AA�����n;�s$�A*�1�����ma�u�\��2�_h%N">�QA��ڈV��1*0�`̌�U���b����=�6A:&�$l����)I�=�|t�p����bcHE'dm�p�	v4�z?���.���"R�����C��!)���Ұf���Ÿ"r���0����cwHޤs8P�.��}�S��nn��|M�E�&�������c�ma]܂�g�cQ����k��1o�P���<%��u'�&n5��ď,d�#f���d�P�X�3��Y���'�JV���B$�({f"Y���Y�rT�2����}���t��b�	�Km/�4p�W�1�����n:K���J�tG���S,l(�V�Z��2�+�@��#*��{�y~ڨ�g�:�+��+���"��d�:�j�U��.y*�^x.�����[L��&}�A��&����
(�ژ3��uW��Z*}g]II;�!�t[��'�za�۶�)����r0QnA��Dܨ�Ԅ�V�/�8J��gpev+.kb*��F�c�:U�d$��m]G��O���JP�\�Xh��џה�� ���?���5�fU7Ȳ[\F3���9���?(ۺ�t�Xv)&сL�ߵ���׵�X\t+��-}�׬�_�Ck�i%/�W�ˬ�a��|KR������겷/V�����"�X��GJ�5'0��¤K�������GfMm0��*���q��z��7�Q��dӣ2��J�Ԉ >b��qi:�>��  �u�d�~�z�E��ѽ�ru^A������&�f��Òv&G��
��4�- ��{u�~����b))�,�;�f�P<�NC�^�������e�<h�W�7ҕ"���$�NBu���BO}�Y�;Q<�Y,�@ >�_� ��#���3C@A9����,����nI>7�m� �b���C�_�il�9�k��r;��躜�=���{�A���(�����G����g.~�ʦ�v^`��V�3�}�!iѽ�%8��x�,ȼ���{V��g�:�+[q1�8��2.�7reo�,���A��N>Zhg:�<�`��}�Ҕx0�F?68�)M��O}����Fr�~�
�o�F��7jGe�G�ӛz��P�@��#����\Z��'������;͏ Eᑸ�v��s�T+]#**����x����c�X�|��zy�	=[z�,�K	�fZ�����p��#~Xh�->B�3���J�h�pu�X���N���l@UG8/�izO	��u�|��[{ov����{��pAʣ�����l}�I�q���ޅX��ib'Ҁ�� u�R�sK�d@� ���O3�G���J���I���Ǵ0m��뇧��Y��N��^����,=�h�zU�tt��jZ%֧mCu�)��[��(ֽH�ʏ{T���3h�o}��0��lb��W:���u��̵�M����$H�P3r�h������ ��R)pF2�;R�썑�J�*�s�Ƿ�U�=�����1pS��WX�21�rq�Ę����q �b|���duk��R�Ex����u��"Bq��?��F�~����d�,�S�&�j�� �;$��(���n�ؗ�1H5����e�Se�n�m�y�l��Ҝ�//`����u��y�&h�'��f'��>*���/KXN���՘�*������K��P^��w�4,l��x�I��$қq�L	��/�?%������*���g}�9f��A��lE���}��K�񠸔�PA���KV����J�l�4��9y��2��2�Tt��u�3�^Lc�f�´�<���u	ש��W���b����K�C*i����u�?M)(y�&�|@}�@�㌊p��;/��S-�`dś�}��rn���i�$M��0�	YcV�)������cnû�gl�L�v�] le���^�Qh�0�/��M�.��ҿ_��P���4O�T��NG\}q?V��v�0o���ep�0Q"\�a��2�жE�oɩ�'�QE���=����u'�TCcݲ�#��A��19�r�0��|�"��rU��@3)���6��ڇ�k��u[J7�Y�ݬ���{R��z2��gO��q�	|̮���ٗѰ<�2�˫A�ح�P�ӆ��}]��y�<�MNDU鼋#�܋%ϫRtpI��W?*Z�
s�Tz�ḥ\���6L��. �i�& A������B0����?�PF��;-�{桔"�c��Tv�-��zRB�W)�F�z(�����?�Q%��M�\����>��ޤ՘��Y�T��:���ل���V�a٤�Q�Z�h+{/b8� 5t��$�+͟�8�+�>������HQ�B`u
���0`�uAs.����f��4�o�V&�i��$"^�6>��-�t��6 pc'�|?�0��v5)���$��U�?�P����,U��Du�&�*�:���"LT�q�,N·�/��`!�Zύ�a���;���8��) ��g��Ĉ�wk����P���a}F��6��0��|�zN;E:��j�@�>p����C7�[��0���`��'��ad�;��3>���o6��|�P�e:�uk��Bɍ5�B&<�߿����R�AJ�߿}[^fM�A���L�嗥̻�ON�W򞌎D�?�R�Jk�:70+?~� �)@���M<�r�b���ՄS��g�#>�ߚ�S�ø��:֝�����Ac2�3z0~A��oO*��Ftכ��X1(#,	a��r�:鋟��~�u�z�B.5k�㋚E��&�B�����#Z�K(�qzf�R�XD�'a٘`���J�1#��ęG>Y6�2g��ft.o�a�U�+�ecu�)I�d�j�k�}�yve�)>��>�~��^/�^��hm���y�h��H�6|ۿ�Ø���&��颌Q�����Xo�!����W��0��+ps�[c߂{zl_�W]���3�AɟoNf�S���9q�y�J$"����p��<�A��~���ғx��J�V$�.]���
@��L����u!#��|���
V��� ?T[�٠KG��/�lZMu�_�A��ӃԱQ1�	�,�5�n��i��0���r�~'Zf�-�W�e�N�j�\D�cU�=�6Ec�'ז�Bz�P4��u��c���?#�u='&��)�����v�P)߸�c�~�2|O{�z�G6IE'>�M�jB�"Φ(�˙AYm@�Z\r/�j`D��/<�m!�`��@>4����n6>��V`/(�%��ޡ����-frPM��J��&՞l�.	����[�ܠ"��=���7��7�A�����h�rꇷ���t}�7-�x[�������O�U��r�J(��d9�t3a�b�[=HQMV�I�!�����_����nꜷ���]e�K���T��A�� �Unc�4��>�`{)�Phco-��s�IH1R����oΑ�7�bi��k~���C����j'9p�v�f^�,-���:�iM(�F���3y�h1�W!����o��S�!�����z�t��6�#���P�ЅO�<��*�N�`^u 1��x���S��sD�p�k���5'}Cj/�RzĲzr��,��܅� ���ŧb��춤$�F�J=��Z�q��8۴�Ib,U�0~�b�#��:U����&���M�L��
��u]��Z��Y�!�A��	�NxolA9���-��0>�9_��'�<�Ȩ"�Y1&(6D�����q�F@Kk�E���f��1JH��M^��2��;����q�xސ�FA�a�q*|rET�����C���C���ӈM�I��Cн\u~���m���{X�$�4o���o���dI�o##�%yy?�W�#��;�ov�0��Λs���'FI�Q��$��B�����m~��q�H��4�m�.U8��!!٧dp�%j�V��g��3?�&
s<�|���F(�;���5�_�RX�_5�=Y]��܎`�'����"�
�$���Y �,����hߠ��Z�Q����S���b:���s爞��D�d��Z�Ƭ?�(�!�RVu����ܪJ�܆�
 ���`��i�Ncꋕ�|�g���F3�iu����0�sy��1����a�`ƹ;�2��y��Ǖ/	?Q���u#Tl���,���%B��ӟ�����ȑ�TVk y��/��i�����^�W��bǅq��m̨��v��c���+<}l�D;��{����d����V��/eF�ec5�o%8yC[��j�^�gy��s�����Ӈye���~G_���˘���~3�}IC>��s��V����O�]�Yg�]�VkJ�����:�� ����"��F��������"��|g��_��&r
,`oc�fL6;�abc��}�n��~,_:ZF��X%�3ΘVٗ�om���cg'(�nx��  j7�2>:�iC�7�K��G�Q$p=�����\��D|O�7h㋮e�Tr��0�"`�s�xI���a�@���sUO�v�O�!=�����'G�5�PM�o�n]:ITԾ��@ �{fȟ�S�o
j�V�[2ߺ���i:�e��!Ze|:6�7M���(��ß���Pg,�D�{����-�ؠ��ac����q����=���PV�����7���IB�Xc҇�ˢ;���J ��ޡm��-kp��L��a�~1���D?����e�C�#M�]���fҟ-�����/�_I��쑂M���q�{��w�w9:%U7lG
�/�?Cӣ�K�:�t������/�F�V���9X4X�g/2�#�%G����m3I�Z2;�iz cr�]�ߚm�X��璮K\��n�wm��*ړ:J�������6BS�\���K��e�0�v旭�Z�U�:=�7��lU���g�;k쳶��e���5�[�G��|�QہL!��5���
��ap~dp����\W����{��皚M<jy}R~�;����3��!|_<g���TsL��T҆��w�ni�?KY/�F����rV m���:ӏ���P.�˷�{����B�>=��9��F�(�5^M��T�B(,�0�3#�|��,�OH��� "w��ِ���8��~��d�j��M�g�w��&`؉E�w��q��I�8��������@F?��O�g|b;�ׇNů��CAda��t8WYv� �4�l�lz�"F�,H�80q�X���v�|ϋb�ڰ��Z���� �7�5q@J�vOf1n��d�m�@
C���K]h��,C��RDz�~�+G�]?���(�'&YE��U�~{c�m�~s�w��ք����*_{?{��lI$���C
���d���l9n>���׈�I������ �M�.��+9��QaMI]�`�Q�93�ro�;�ݝ����c	���Db��OAԌ*g?A轘���ѧ/�v� 8��ؼ�B}<�LAo�9�D_n�5�`!_��u�Wi���ajZ|�&��Z�#�)/v��h�������Cńl�8b�X:�f���F�8߶cF�#a�,n���.	l<q4d�$ȇ��\b�#�1Q�	�v*jRL����ӆ'�<h@�*�g<Z��X�(�P�Usˣ�f��P����P�>y5<�B�?"�Τ�1�]���n�M��T�S/d[��⹼����y��"z^�h�x\��j��_J؃yn����(	����6$Ad���T~{��.�^Vw���#�gΑ��>�ى������rU�:'jb��)RNܹ	*&�O��vC�8�Փ%��$�g���!�!u� �X��۬�u�eup+V�������^�C�j��Gݷ��#�dIC�I�kߘ��bz-
=Sd���ƥ���͇��h�ACb��c�����DXXՕXӘ�%��8��f.���I�j-�(R�&�8�l��ᬍN�r1)U�!�:��2�y�T����{>o�b���s�c*�cu�������／����CՉF��pE�����6���o��o��Q>+	j�Z$7k���i���6� ��1|ܓ�7�fl2�3���C���,�`��Z{�r�<mI�
�e��Ց)ն��]���S�$��]�eT��}���:�aS r6���f�����D�^��?1G%r��.�I�?�����t�y�;��\��\@?b/��}��>��*����8��P���g��w��Y�"� �1^�Y�ޞݼ�	����H��pa�ד����' Ľ"4dm�UF�v����	���Hlڌ\ؚ+��
$��m^���G�4ֵ�����Vx2%JdV�>�p���Tҕ�K6׎.���r?��rZ�D]���T�a|���{7����$	�	�%fN�˥@3�c���+#���`���,�@\D-�$`w?!���݆E����>����V�Rҋe�N�Rk�#�ٺ���k/��0{�
̪��W�P)7�M�[��oγym�7�/����ݎ&?��,"�P��w~�݉�*����jA��\g��nuZfV����3J^�l�)�\@P�*MÎ�v%��&04^��;x����R���O��:I0G�KL��zG��P��1N�>Duԣ�t>�-�&Us������e(����y����qT0>����S��R�ĔiN��~�c��H���[�@~��j&c��ڨ{rL1�B�����?���hJ�b[a� �s"%�Z
�a��.�E�Hlބ��/� Q	�&Kq�Β�9%1x� 9c���ײ����!�N>�;���n{C+�9cx��i�o�e�+���BO�&OS�z׼D'��x,vy�,)��ڦW��4�&2��e)�Ny���4=���J%�h�h�Ji��i�ibY��jMܽ�\��[J+���ڥH�p\���ț��o�_�`^ZL�ڿ!QW�I�u�H���̩��mZ�����+�|�+<���χ>LuT_���"�}�^xI�x�ྜ��(r�y�k���#��
���ڡ@{�w�*��0�C��t^s�<��$S�����D��r�Bd8k��������%�����Q4�?������E���s`ŭ�	q������6�sy�����*g2^[n�QM���p]l|�����ꡦ�oC������¾k���G�!���k=�VMK���#x�)x����A�����n�P)���tO�F^�8��ۚ=|�����~b�'�?�o�����H±�D-�&Iz���|�7!a%�j��( ~����=����bA}I�����Z�2;{%��kb�����S��RF��C!Z���&� �xy�J%�F�ԫ��:Meш'�"c[$�w��M�e�.���#@�泱��G�q�)�R�x	�G=���_1myxr��s��"0���"�"S��Gy"�B�]�Q\�׼*�ο0,�W˨�?)��}dV��kh�E+>�K(�]���:t�ط��B�4�߲B�!e&K/���`F��q���t�=�����o�/f��=>��C�c����U�i�p�
����o����W�ǎ<.&���s�H�dHYX+}�/
�E(2�5��_VʼZ�^p����R���SO�*v�o"���Z��|�3H�F���>Ȏļ��D�xX�����,� ����-|H��"8��X�Z��B�Cs�u��i:H!��B������^��)0&JV�a�M�FK���j���{l5��:�T�����Q�P�cұWm����./ZћZ1 ��|�y+�@#-֏;�{��gK/�kT�=h���C{��2N��9�5H�h=F|��K����qO!��	{�P&����7���'r��H:�2�s�����P9/4\��B��z��~b1���ɝZ�cK�ݵ��a�w�[���B�ꝷ�ʆ�59M�R{��y��G#��J�.�C��x�fA�ʗ�\w���[\U�xw�F�l�3����?>�%�m�s���EŇ���B�8y�����B6)��.N&�����4�Zz�V�P�����W-���O�J�8ÄVD���R�Wہ����+4۴Yx���f����I�IÁka�2�z�����B������0`��C�}��e��q�@�:X�T���ɦ�I(Il���Ј)zh��z�I�"���b�:fѧҞ"��Jz��Q@X���E���l�6N�a`IU�t�A����k�T��q>DV+��N(yr�b^S�|
��QG��g܁$�c��Q��&0�* G���W�j�h�Or�͢�>ҙ���O�W=��M�"�
�An5M�HfK�ߜ�Eu������L�,�! �R�\0p�g�7��N[i�A�B2�f��˼�dU�?��`�-<B���,X>*C���K�{��W=��"���%���[pn�N���[��� Q�D#>�<��=�G ND:�r��76���M��B3��ʸO w©�L�����TŅ��h��<�@�G�]!��ާ�^E���tq <���B�\{h��0.�3�����C�֣��΋B��<���i��Y�]�,[�QQ���N6���t�L�2��#� �pRTbi?1S����KAW�5�����6A���%�����	����;�����h\*�Ou�±��yj�>�y`�ЕI�Na3d��vW�)�:��@��:?�F԰0���%�8_���Lk�r��os~}W�ᡢW�\���xkm���⎰hX���`j�&O*�!BD�H��3���N� ����X� �ƿP\ۥ���P��R�jb�>��J֎���E���>S �Uy�jMg��0�c�N� �6�@x��~(he͙�]d{+�n�D��N6�����^BӮXU���DY:�(A^��V�CȮb�?�i'#��u�NľpmqF�J@.�qpK@=�r��j�Kå|nޣ����)0���Cssɢ(�q�+�΄�qYъ��6�++u~���Z����	���c�w���-�OA8�,&����)e}�W]��o�[�t���7�$�5<���+�O\�w�`o�S)�J+iC�[�gs�;��I�aE��Q��Pj�
j#�u�=�(tIV,'�э�C_�Q7؋��J?�6}���~��L;�9c�1�r]s��~����q�emîu d"l���B(�s>X��a��=�0���7 ,#w=����r����6��S�C �ʺ�_<����{��,��e�ہ�d��]��}���"�Z����H��,:�x�zսF�Ӏ�Z������/����n��1�Rϧz��Sܷ������)C�
J)���:,+�%�D��4�e��=��y\���v�s@�6��S��*B�b��`�cU����9f�����u�^�A�OЦ��"��Y��������?���1�j��@ɑ"a�p}�*2����/9�l��M>��5m�5�^�w��	(r�N���PK�����) td�2�A`� �5�@�eP�_�]�ۊr:��>.�X�Z��� �H�N� ��P3�a� ����9H/����*�4c�#r��@p���8j�D-Ç�yMMU�ۓs���7aՅ�!ꚪ{���tuZ��i����E��\D	���r�O����S�C]�D/��P�f�T��>��s��ܓ��m�)q̿�O�8��T�P`��%ŭK)J��dJ�gy����E6�eg�	!C.i�Õ
&�δ�g�K��o�$v I��d4�.	DY�Uf'���m�̎fPt&b�����us�x�!�z�����5�7*4��g����=��OC�X���+�7�g��~+����M��H;�Ġ7��=�=�G'�˵J��^u}��� ���1�r�K �@�'6�<���yY�
�I;��/�6�,�UZ�GV=����ѧ�����pLOú{�*W!�������}��Υ��¡P�݀ۺ����+��h��z��[�W��b1Ē(k�W\Dq�M�|:�R�Zz�Ym�����[� |ƣ��!9�9j�p�fEX�ؘ4i����::yV��ӧZjvR����b�8�H�f!���qJ�*�94���
P� 	U����	X��|l���Qp2!9�,W��u�pU�n[��UՖ�<$҇ ��̖zT�rH�r�!�w�j�h�ٽ���?������,8��	�|��i���J 32���B�a���D7�,C!�ÑLv��}2`.��e�{W\3��G�MeiB���lNb�9�nX�YuǾ�����%�d�����t�7��B�z��}���wl=��MG�p,���$�ux<��ÀQ���Z��ٳ2�쁢.w\7y�M�t�0�/���nǶMVH:X��FƗGJ�"��;�s'�\��?^z�Y�$�NC�}�F�|FP�`��P�^�&�˰��5-E/V�_d>-pqI��M�3�+��;�W�=�ȱ&�T�a0b����S�=�ދW��9��;Ԅ_��*�D�uBw�v*�G5<E��;	˾���֡w�v��G�ץ#z�^�t�-�F$4�NS#DEb�`m�6��h���ϼ@h��;�!2ڐ"�uUۃy�Si�p���O/рt\��n�Xh�l7Љ�H^���[��C�=�JnT��H��ф���+��x@�ԧ?�!s`͏���q�=f.ͷ+�8y��Q�]F����!r�Š��M�~֦ !՜�}#�#pg���{���y3d�[�2-�\ /~�v�5VQ������8�o�
JV���\�>�Ǜ ����d�C���_\��٢y���7�^Og����P��>���	V
����Ǌ�@���q3=��H<!i����>��\�ү�^u\����ّ1K��h�gO7����WH��/�1^Y<�{�b(���1p�k�����}�ņ
&K&ԟ (��L5t���4ި�n[V�*4�l��漑�$�[�B�SI��y,3�'Oh��;�&�mu�2��}�;�%)S����0����d&5'�Ы]	�Q^tW��b)���ũ��C26���<�烱�0{�"E��1t�	���t��tU���F�x"7���Z^�1>�3�Qm,(TV�	��ɭrx|�;?)µ�-�:b�./m,��DQ^����wŤ��S����(�)�0,KX�ϵ�@Z� ��s��F�M��U^#$[���v7N@�|�S��cP}j^���,-���N�";>�J�\1O�����(e`Wp�[a��c�̡��5l��~���Z�`Bl�$��^}��Z�ƌ%�ѡg��{��D(�T�?^���ە����^��omO[G�v�N���v��ӻ�	dw��3W:nt���z"���A�2C����nh^���Ά�,���5�}�j������һ��[6*����T�|���bU�#E�D���s�7���pV��].�]���>fǽ����q���UG�9�Of�Ͻ�*@ui%Ett6���д1�l�9��4�cv��^][���ԋ�]'�oܭ�wL��T��q|�Òn��Au_��(i�	4�c����ʑN0Dm-Md=s�9P���3��j_�$��ef�Lľ��idP���i�c޸R�����U\u3�	�_��>ĳS���T+�˩[�R색O�8<�b����]�kg?qD�z�lؗ�Z�ꀽ_�6>O�S���3O.�r����C;��Z���.�>���,�Ĥq��p�}�X\�����i�D�0t�x@��P�!Xq��&i�E�.�v�!=沢ɾ@L��l�*�S���t�X�G&P'�f�P��8Z�|�.�X�B?���{�${�������H���!����۶,�Y��H�S]��vԏ�[��(E�ݕ\8pV�g�!2D#S�fU͞UN/f4����
�ƥ����P�ĉ�%�F����S.��z$��V�ݢ<[������7&�(~[��<$���UN���B`�D/]=^�B57�Q��ɲ��r�	��|���F�|:��̱ �M���3-?�����jjH{��Z�f��[�5`��_2����g3B���H�E��9�q�f2�(�7@ܬ�f��h7��p��8�|;|��^Xv"D;kh�$,�G�F��*�� ����g���t��jێ�࿐�0�m�_r�3&D�Ӟ
_"j݊;�<��0�A�{�}�LW�>�X(=�E�2�ذġ�cګ3r�)���y,�',�"�.�����u��c��������J?�~���I�9ka�P���DT����[���@!�����5�8*[x�AV��,
(
o7�X�$g�&A��������R�k�����T�Q' @��G>괲������/�T(��x��P��Qp�u)������	b��e�D|��}_��Y��Ъ���{H���Fb)� v���xFң�_�+�%i.:�v�p�[ ���\4[��ؚ(F#�c�8e���*��e�0��c8�@��|����&����E�ܛ3��:���V���m!e(�ށ�vӕW�o����Q�%[N�و����E�Ĉo®>�x��5��Ɨ,'���`[C�ǁB�)܅�7��\��c�I��v?Y�������zZ)�d"�/� �xs��0W�Q,�/�U�T|Rf�w�Z�����Q;����� [y�鉊�[f�J�ov���ūy_��u����wj2�BK��g3�
`�_n]~+�`������G9V#&���Mw5v�g'*�;�8��֭TI�}6H�(�ـ+l�W�5�>1�Iy
]ذ�Cc v����y�{��P��>a�J��9��s�^�'�>u��ZA���z�E(c�e='�-e�+��O�h��B�z�o��7�0x�\��wg��bB����9��1'�b��BA�<<	��_&�)NYR�햣.�Hb8��4b�U b�����%�-7�;1�Mǅ �߀�z����Ѳ�X�nݴ�b!� �cCW���C�u$I�K��\�,��GO*�l3����&�P�y������+���8˫�_�i�?�3�%]Y��qPY�6 ��{"j����?��eY�3+������ TS;�Yu4V�
����m�7�w߽߷4�-��
ڽ��z��y0	@Ԥ�*S6��A����bt��o��7��(\�&_�_�[���\��g����ݦ�H�)�H�c	�S�d�7��"�=��Sw���&�������K��p�R��djUX�n�̀��O�B�	G_Z����ki�7���	�j��9�I�-���4В��l�E�j<��
lM�9�)�1��(a-�`�m����B����{{M���g=+9T`UƦ��A�j��3�l��A�.ݹ������r������7�A��ɉ%����#AП�$��[3��N(t� E�t��C��-N����������s{��Is����]I�5�f�
/hp� �a*���}��G�*�s#C~�_[��Hexἇ�1�E�[]�����X8�1�!��5
O���׾*e䶼d��H*M �3Q���;�h�7�=�{�=��U�?����<�ϗF4�&��̻�hz���e���tQ�J��$�Z�u���gu՝�t/�uw�F���ŮƤ3�\x{m㙆�\���3�1)��ڃ���m�L ��ȴ�,iF,�@�0����$�<�Y|�~�tu_N�Wg5�MkTަ}�j ����ۂr����)Jҗp��ǁ#\B�U��z&��X�����4�~<�'g"֬׸w�l�{�V�l���/��͆\Ld@�Y�pߎ1���d�����wM�Vǥ8�f$��)A��G{�������z\�����k>��M�E��yM;��`��Tns2*LCEx�-?�]��K��y�hR��}����ׯ�8Y����챀,ӹ���əZ�K�J*�3�!.I�J5�S}�� W�����5�4B��?6W�t1ƌMc�Gz���H�@����
���@�=}��k%n���cW�{��yL�'K���v�~T&4��Vl�ᑌ���̇v�ZOQ�!b��z�X7�4bt+IK�Z��9
T�(����	Q��9
u@��⍩�X�Fsb%Ȏ-�W���<����9W�X�$S؂�B�ь�8�y˾�X'��L���Ϧ1���"�5!�)_)����y���>,Z����p;����o�gC�*��p7@�:��j5$�()�@Um������=vR���-�4@�e+kڄ�W6ؽs��>�,�(�U� `}����u��1�\��[��82["�J������@[���|��ii�WmvM�t�9�X\���lE��U�Y��,�t'� ���>8v.�E԰'k�8�]?K7=�3C�$�&^9x�68���lq��2�N��շ|�c����y�� �㭝Lt ,�{z�!�ʰ�pj����zR"�@|I��b%�!1�f�Ꙛ+�x )a۴� ;�3?�0+7-���(�+�e���^>�ാ�2ϝ�C+����X����n=����a`PrJZB�h�n���e�O����>=�q ���P����Ñ3$���
�87���)N��bE�I=� ��7�o����Y�tZ�䤓��_V��u�I>P�D����o7��I��{��-���;��)믗�k0�G>�*�<�7Eu��#���}䄶
Q
�&J"�ǧ�ÿ�i:��H���O��m�%ao�;�<G�4�^3u��������}��*-��3��û�=3��ZpGX�??:
լ���!�� ��m(��M�9H�1eՀ�CA`j�m1G�!���iRq�ms�����F*��Ef�{5$	�d�ԡ_!V ���:=O�����©&/p��:�S2>�����ˌ��4	?ͬ��N��*���S\ ��F�(��dD��.(����U}eW��V*YX�t�	�(+]�+r�j<��6�ڪ���)����Ϟ,� �{����c���q�C��D{jW�o_?y�6ja`cc�E�}C`�^�YX���T�߇�i)��ݨ�#��m��Yy�8n�CA�0��y�>Gd��\)����]*�3+����K3��8����a����no�܆�"�җ��Z���,���l�J����;��aN���< ��1�W��)�+g] �,��4^Ͱ��Gk<��$�M'M�P;���}^�ׇY��}�b�L	.J���k=���o�1ڵ*ğ�5F`bV���#�2U���@^�����GѴq@�͍A�¿��=�u��RY�)�w�Em�x���1��n�4-B�Zk}���d���ryU�D�6[�I�
�ae��*�`W/�t|��	z!X��d�g���G�5���ic��1�=kL��b'���ɤ#��VG(;�7�}��os�\h�@y� C���h�t'F�f��Ĥ���q��J��4�O*�A�C��E�T�����8��~$QE���V���/�?3�����Oa�}���3j�K��g���g���7n��������c"��if<�nIj�nS��t(��G��Xw�4�u��B^4n1�k�ZQ����W��j�w��-�Y�qc�
WC�qH����̢en����jK���|���0ծ����[����PN'r�hy�͌!H���������G�q�&LMГ��L�ַLJ�TAs�RT���OL�A��,a�¨ X^#A�{n�5G��Uc�O�?7�Kx�����ﻑ.�<e43���QF5����0�G�M���U�o v�(�xg6m��C�mՒ�C�`W,�-�Z
e�i�{�]3l�⸞���19��M��6E�o�7���"9E9��O���������$��Rʮ�䪗t��f�p�{��[Dɲ@��^�$���d���aT�L�5pp�[��]D�3��Q��`YJ�#?�@����G���r6���I������SU/<A��3Y{!�|�a}��Ӕǩ:�%q||WqH�`q��rW�<W���YF��M�g:Ȱ\.|��]�����8,9��qs<B�i���_��"�s��]M�$�=B���0�\#dV1�Ͽ�-�|�Aodj�g*�a%�f0k6�S}s����Pg}�@lE��5��?��I�dUV|�1mL�]�`q=�>���Z,.�E�7��?d���E��V@�?V��ӿ�0
r6$�%�/)��i���b��+i��lK�6a@�p'��04i�=S�{�Uf.w�2�R���7�� ��!��'�s�Ԓ~�l�;���ĽS+t/�{�Ђ���8��@6�S�%R����m��r���~�א�
�2Yp���
� \t�It[L����ї��}6����i����$F��)vwZ��1�8a��")�`]�LE���X �à�dy�!Z��?�(�R���C&B�\��g�WB�C&�2YF;%0&��x} 5�����8�M�l~�������V>l;�������]�`�[Ų�J�,]~"��oP��4��%�Il��x�������	#wn`X��a�
���E�K�/����;�a~��k@5�!��J���l�l�����Z]+T���9x�,�t�t ��.�G��h?�1$|��r���FQ��(�ƶ9��ђ�J���5�,���s]_�t����`c���DI��ĝ��f8Sc�N<4�gs�4�$o��E�$�>/�	w`�+ˇu�C���_�vR�0l�Y�-�B�K��ȝ��%-v]b~?����~�!��p��!л�W���xz(�ل����F�83�?���%���:�P�Z���������l�#:羽z���9��8a��Z�5+y��.����V��k� ���n�c���>nw�������+��c���G9��pjzЯ�(���?5�\fGm�y��{�(uFci�.��� ���'H��ҟ��8�U-��	$�i��6A-��I�^p<t���m�r�w �l��%R���ܛ{I��oL������k}G�+����9��e��*^���2M��YK�� �`��`|�.�ᢦ�{#[2[:�Y�)��8�2�S��L���+��K_�]^Éf?�`-R���5WZx����*o�z�GPg����e�#H	�V����J�/<��(���z�4<Tl��@eg~z��-,��ʩY�'k�5�4���t�zz�*wQk[0qJ�J�;>�5E���Y�0�K���ys�9�N�oڼ�����=HnU�q_ےk�-�א��M���8���<�����x�g(R��>�E���W��@m��N7
����J� ��Ǚ(����[�0�u�[Έ��E�m���nC��f��b!␿�Qۇ�p��R�ɤ�s���ޠ�݂�N(J���E�[��J�r�[�`E\-�*}u��Q�9*�Sh�b Ll�s���"o��EX�#=ՉS��^"��/�Ee��Z"�+=�9��䋤�\�R�·Gȫ0*G������"����%��~D���ԧ�������<���N#�G�^��8P�'�W�k���6�)'�$l��Iq�22���N�>���� $��r.��E���Y�|�k	�G��[�*�0}e�m�Y�'��n��/^��k.:k�.Ԗ��pI�;��lX�9�1�4�{��$�i�!��@�=�,�Nhr�5S���N����� ��|*�B���J�u�����l6`B��DH���QO:�볷��:�]�}�w�?�v��������P\���[�B9����c���)�+�0�-���'�5��O�]Rj�oY�<iϡIr�mՇ<��T�L�B�������F$ɖ�_��3P*Ͼ\k�����;	�T4}�n�~Xm��%9UaI�Ԥ�wVq�&��������zl�Uû����K���{��nTon��gD��{u�2��,�0�f���I1��$5�vO�-�YB��p%6~��m˝@V�8�<��!_R�gMGh� J��)��w�5D�k:��6?��<K�����r��j1 �
J�_NG̙p�@ml�@5"tGs&�9@��� ÿ�����x9�9.������`J��\x�:�X� �H�0�<�gXq~"��F��R�|�����������g�KR�*�i��o���� ��*_!}�n�/V:Kn��!��$h.C]���
�j  �+ˀMA(᏿��/���Ņ��nƆ��֪):�v�Y/35(�z�rkR=���brnYH.�Ĩ\�]��	6`=��Pn� �(����.��˵���Bx��v�Gt-Hx��(�;;������}�}�rؖ*�/8��	��8���1�N{|"��A�^��T����-���kc�ɱ~�{?�vT�rJvחd�:���]����3��6s�

���H��J�m�|4����s��Z��	<M)��g��[�+��F�#v��"XM��k�j�04C8�دsj3�|� �|B�]�m��ēE�\�|�J�v��"`w�s���봘-8q�eo���-�*�4�<iP�"#*��*�:z��6
�9P�S�	�f�}:�Cz��������1��}������ts��+7�������UJ瓁��� w����J�ئ����|�Vit7����`����j�q�4d�RI�����<
y�oz*���au�wK������	\y�Å�*Ǔ��͋��OՀ�	���*���o� �9罓�[��[c2�H��iU�]5;�J.Ƭ�y@:�du�^�z
�Y��0��ٙ�,B�A����0�!�f	˶S��=G��^ul	8�q>���/���q�BÆ"���_HlwB��S^0��:�Ú
����r !@���@A,7�}{v����.�/20�lQQ��*��]~� �7vK�@s��]���L�y�E f�F�7��U*l�Ze��sΌ\�ߢ��$�����e�8�9ed3�w%��қvjptU�}��VӪc���H��n�I���W��mƑ���A��o2�pӌS�@ONА�Fu�Mq�6��2B1��֘:zswl6C:�"�K��������uǧ��w!	G�:��{1ʈA�W$>YCc���]�~�9�`!���|r ;֣�������Àt�r��^��l&Ym��[䚟U���R��&�09@t�����I9����r���{�A	ǹ��7*�d��{�����$Tם�o��Mu� ��5�C�jW�o�&uէó�5S<��k�}���Ƃ6Ґ
�a��+��ë�db�%:��{�F͢�?�|9A�Ծh�ru-�!�f[��:�����,�)+���@���V㞉}�t)�__�O�������i��Ω�g޲?�#I�w��<L\�nҡK2xí+�>Q:�cͲ�L��+Ȑ�(�L�\b��?�:��s�z���Oab`��N!'G�Fc4q� Z��y4�:��GÔ̄�s���m�!���C��(�/���5n��N�m���[E�O�����9y6��55�Z"���&SM��)4bm��V[j�!KKs�P	���U�D]oPF��I<�@��Ǭ�eR�k$��yB����
������粱�e�2���-)���)��ˋT8�M��C���(� i:+���Y"vpm�v´����h��3�� �T8� ���b��ə����`cЎ����=��`�hp�H����|S�C�Eb}��M�-������NC�x��l_w���i��VP�u7/*��Qk�rp�O�l
� j^����j��� 3|ِ7K��f��}&�RBN��"1�,�r����m�X{n�ݰKP�4-��1�ݛ�r��rS)U�� zn�A�CK��_4r�`�[һ%��s�I̤�s`5�w>���g�<lUٸn�f~�$7!�Cu���\B�����sTf��,��w����;�>���w!�&AǼH���4���������S���])#��_����uX�*H��aj�C���v�6�n��]H�Rc_�{?�E�T�������K�0��'k!���@'-iI�5W��󤇮��k?n���6�н!�
j�_
��N���6����	�����m��uD0���hbW�]k�.�h�O刀F�,��hs�5Ds���CvML�Q�qR�`��_�LL�1�x�C����-X��*�k_ҩ|eT�#���'.�/�Y��zD��d'O��&@�#!O+2v��%���=<�M�]Ź;�Ys�0��.lY�TD>HNG�AdI���0A�w(�p.%�"4��a�C�T�R�M���*�)�}zÝ�d��c�hl�j���Z[@.ו���C��8~0>�9���T�t�n�ry�t�2�E"9�fN?�#��t����F�,6J�BU��#E��L�fK���͐�c7�J�˩�ƙ⤃�wj�Ե��Ȃv�f�T�>e��ru9A�e��N>2�*����)>[���b�-evE`���q�3X��:��;g��}�3� /ƱH/�F�����~'�Y�bA�Ƞc���(��R���� ǲ8qĻn.�Ua�j>�ႝ
�$�U�h�	Q|��7Q{Z�/LΤq����Ҁ�R-OT�5�h+��T���]���uC�t���qǃJ8׳R���ip>`��G�x��RS�[�I�� e=o�%	�2����	�o_����m@#��L�G~���S��{���DDĢk�)R[C�#���O2i�a���{(^�	w���h+j[��hգ[2��3�O�s��a�
��k�s��m�ǘy�59}��Na).e=g���N;��y(�8�}���G�lV��B��K�g*�t��!4��谷\;ۏ|u߇�Z�j 71��B�Y���0Ȗ���s�̜�X ���N����1�����\�W�RtZ��~�g�R-1s˙�z�1�a���UV�\{j`������ (�
VK�V����Q��Pt�q^e�Y��	3��9�Jw�n��A��'��o��v�� �w����Z"��"�|�_�
1�p H�n�V;�w����6��kx?�Rs\�덇z���΁�{��b�bb!�Az�q��D09C��P�C:�q�.LZS�Q~G���Y�!�:����ߚ%��o8%��s�B��m�z�v����������iTp(��c�x��`�V�fH$w��wz���� �.B��ᶵ�bd��s�BzgyM��Bᜀ��d�9�E���(Mzۋ���h	��Vo��X#�*�b�L�p[��=u����H>"�?�)��l����S�s�����1�0�V��ؓ��Qgoý(b&��Mf� ��b�@��&�TR��=9ǰ�>�Ւ�	IMh�p�<o��cGv�'�Ɓ�?�$�XW��P�!�4���Y�VA����DO�����.hn���V6@⎢i��� ~�^��)ʗ��Hg�vM�w��چ��n�n�O`C��`q����[��rkD#0��O3����u����� ��*/a[���Ms�9.���Uu���.� ���:e3'���j��%�E⥧������K��FV b���u����1Ĩ3�s�jȧ;�]-�q��`�;�oQz�mG�8vi��M�CC�	Q��k%H���j�ǽ܃|�����&bM����DAe�%���t�����)RV��1��jRU�AUB!FEL�-���I)�^^��[n>�,��*wp8���y�������Y��O�^�o�t;�;(�i�K� � *#�:�='�luOi�~W������L��[ܽ�F�{�ֲ~x�yL��uÇ�b�$�	��\DN[zβ���!�yOEb�|�DT'zl�!2�\ ��3!�v�V�`�o�!�ˑc�e*j���o�.%$&�|�I�JKp{w�(+6���o�(~j��9��fw"��`N�~��g�����ڊt�A$pAg
:颥Y�57�5��	7`�>gh�k5�:�� ��W�\����NΙ��W�0E���9(-%�60/ؾb g7�jY��O|X�{l�� ��u��)Q��ʵ��Vݰ�t2��|�<�厎L�/0=8[c�� *-n�KG�D2�j	5<1!��#���Ea�����o�}s�r�ݮ����Y@�C���,�8�h�{�wB,H�+m{$a��zl ��{nn��rI��kC�J��k��ɇ��3�,��U	D���ü)VMe� כ^�����ρ8���I�d+eqTȴy���C�PB/L���2L������I��(T��GNKW��6����c �ݶ�}t�Kɣ���͕�!��L�@���S�j�|���l���v$��r}+���г����2�`��o�"M�#dQ�/Z�7I̋�%�~]�~jp4�D���]ޒ}t��?���"4�Q5��f݌^�%���p?���)iw^�͝~� L� <';���|�
�;���¶������9���"D�Ħ8ǁr��.�S?=ɔDy������_M�����X8vN��O]�P3�i�3#�_�y�r6�_ѸG-|VV��'�Mٚ a�jY�[2�������ܭ(���[�¥��s��r<d.G��O� �K|���O�/�Y)�.&3|�|��ئ�o��8��/�!�܃��e�F�ı���1��5E[,m��a|������-�S�E�|�H�H����;	w-��MA�޼pp!��	l��%�"�/?��w�ӹ��^`�ᓈ�&-�?"Lc�5��<���A���`��8Δ�sT�0��R�r�<q>$Z�'cr+����?�	���;g���w ��>OA�(��yG�����q
���
���[Fk������3l��M.��5b��1����`����`�ycg�y ����Ւ|O��k(���3$�J(���KU�w�@���"���pX�|Ԯ%�pV}^^������neP�^އH��O�H���U,c�Ͽ���8@1L Ʈ���%����d�,v�;3���*�!�pY��N�����@N|�i��)ɲ���x���G�Ȇ��죄`�f@}�b�ei���J�pM��c��a�_���fTe$�/�!�glxA0{U?��9��l�.�Iv�$����D\�ڟF9L�?�2i�z��#+'ڶq�۷��w�<���s��/�f��3�Mu���+�~�Y�w
�K�(�*��޶ۣ�L�B#��qy }��`l��5C�ba���� U-�Q셯�F�¢I���=�B�V-����Ehd�����@�$�'s���U�����}�c��d����?���6�R"�[�:t�4C���fr���tK��.V+5@\�^ϗ:�"�Ɯ�&U5�����;a��e���/J�<vu�Y�M��Q�;����J��K���uc6���E��UI{����=��+�7(e��T��ݝ����n�A��'�tK�Q�p�����Y�J}'��lu2��c�q�������4QYZ�po�����%�	�~fl�1 Sa�,^�w�������1���l��1m���.�M�UgO� !?j�{�2��Q��O�W�i�K����i�䡕�ļ5?DR��#Ѣ�W.���&B�;�7aprr5ߠ�'A���"	��M�Z�5<l�!�#��RT1цl�$6Y��N�8���G���s�77�M��z����ן�^Ƒ��3J�һz��h{�労	[�7��֝cD�[;Y���F�����G�u`�
��ƈ���G�Kx'�5ՒH�G۩�'����ʊ��Q��E�H����j���֊�!�!��!��7��n���DD.J�]@3�cf
��{���TdPh����z�5��M�(G�s�K*ӗ.�?�Z���_M��XiD8\�P"���^PI�b��:tt��|[�5�c�m�4m����C��Q_fGb��D���L	�����z��"�Co���]ld�M��n�R/���8�f!�;h�w�iӚȾz=�� �;�wN��m�Tt�BC�����2~ҏt����9�k��z!��H.�M2b�Z�eR4�Ц�����I�L���CN����J*W����$�+����꜋}�F��mX�
C�?+��pou�+��^s5�8b�[���l�R�5�������+r�uTA5�Meƅ7�0O߇�8�摍������t`�g��gTٗ���s5����UQ8�b�r�y���=���v��/�G��]B�ݢ��u���H/������U�R0柉3��uD�0�rЎ�1����=�J�My҇��}�]!$�jE��f y���@�������R�<��u��0~'=�z��9��QG[,C\��gu0�T
�i�`���H�T^��^��+G-푞��u��S�O�	{��R�[1D`���Ʌ(�c���'sH˓,z1ǟ����u z� !|�xPc��!����I�����Q,$'�Z��<��qB{���o�Q��H!�x�Z\��
�_����D�@CnCA�S���\27��"�#�ԥ���W&���׍��Ce��YD���m$k����I����Ӷ�#W+�)O���s����&\6X�����>�����H���A;n2���r)�a��ɨ��!P��d�Y�>$-��H�v̊�>�i�}F,���Q�/��<��|:�-����l,�R���%�o;���"C�
������ě�,��N�֘�H�?j���@�M�2~�P� Nr|y��eZ/�
��|���[@^!��JؿW|\��Ӻi"z����M��2����:�����4���:O�c��0��o7"�{s��DI!N��+�#!��g��i�R�d%��]A���6�X=���
	!O���&Rͽ�&P#�%�Q�T���8jDR1�ϫ���e-�[	ŀ2ą&���gR"t��w�]$�4�ڼc�Ɍ�7�r*���OP���5�)��\��ې���G!Fe���(�2�W�{G���Y�.���g�>A��+,�:hr9}���E'7a���+/�5��U��[���%��b1f�n��i��8�2@�Ԡ�5��*2�ȣ�M�x!���1��̈�',��Q�a9�-^�wu�����d�A�s,�󃃇��Tr�Z�ʫC�Z����D�i��]ǻ���B������v9M	9�����#�'�������X����";��y��7Sݎ�����/�Ӱ7�A�M���������� S�2�Y4v���M{����h���~F�a+q@�w�ԋ�l�R(Qc[u��I�*pǫ��@�?��+W��=�}솏����ln4�eO�q8TRʼWSn��iv���>��
Ri���gL"��;�B�&Ӛ'�IP�V�x���g��r��&��c���cF�����$i�D�{f�Ʉ��#Y�R:Ns�	I�����t�^Z�.��z���D	�[���N�����7f]O��#��s�UBQ)mn�8���<�㴬���u��I�3_��/-�M�U�dTC!�T���7}�h��քf�z��f<+�\�R/�p�z�^���yR�&WF��P�Yr�{�eu�>R���YM0k��Mƿ�����} ��K�D�R��5P$EzQ���q'E������[��MJ	��/+�-�1-,O�O���s͡�B���	�]Ac/V�"��:�ST��.�\6	����xP�D���7Rȯ�6s �V)�:m���������gA[|�Q���O�����y�2�G���vH�V�gS�@d�����6@��-f�v7)I��J�Rx{%���Q�K�bX�͊���Ԇ�ÿ��K�(U��}����[qlge��;�Lc�~u
W�뚥:��I�8 jZ��]���?�@e�;�p������}�J�����t��zI"�~�c���L�]��S΀�k�*2��R��V��� ��:�zs̣��>�8�Oer@�"���K�jY��f�]�c�4);�Q0����X�
?���Z���1���æ��2���(YJBFJ�W�Au�;���O0�W{[��$n뉫�L9ٷ�ˬ�-����%����y���* s�O�v�X�@��J� /�����RI�r8[�b^7��&.H�B5�ޠ�8����pko�hH�8�2&���j��gR�u��|��fP�E�p�)�Ņ�=�$]s������F��(�	总�'�\UU�,�����^��'�q���/Y�����г���������}�T�z�R�{9m��Ow���X}RQoI�E��\����@�V�F�����n��'~#t`ua���j+$ˤ��U��1糘��Q��p�)[dOS�o��' .�<�^�l7�����r&P�	��7�c���������:�]&�J%�H��.��4Y���3���D��\7�=���'����A6���Y�t}~}�AQH� ���P��pb�������a��LMo���H��q��Y�5KF*��� �
�6)Q�%�F�3<��;�q(�T�k;'0�T^��Q����d/��3jm�	��E�W�O����v� xǘ+�50}����Z�Hi���x���m���. ��T��A��ex^����m:�����C��(8�d;�5��b�ͳi��%�iN����"��v�O��Rl��qi�]�����Ia�|���]��F�کMF<�)�wׅP��?���p̀$�&4�o�l�EX�zB�݉�;C��D��ГW�c�d��_��{o�` O��F��JaI�;��}����B[���=��K��;��sD|1$� �����"��g���.���MU�8�W�����۲l��C����Vc��y�Ϻ ��e��p�&��W ���2���{-���w5X6��ϧ�f^f��'Q�̄j����n�\�r�ƨ	p�[<}���9AnŠX`!!D*m,�^B��M�M�I��>�`���Q�p�V�Z7����H,��̱���%���DL���֎1�bP������ꚐX~}X�@��\����x�P���J���Y��E���y�3���;V�����^��BF��v%�v�=��if���HKg#A`�2��T�c__;�⮌}Sbw����T��"j�W��G�J�6�Gic9��!�"�3bQ�	�?%sL�8'�Z^��/-��O��7�Sz��hU��-��i"�s�K?y����ǁ*�MV��8��)8��,��p|�����M��G$q�^#i�R,.������K��E����tdd)�z�������� [W|f�(��о �//���7>Uܑ�I�������G?ImL�� ��궳�y����ɨs�,����Q�Z����f��ό_.9b#����,��.�fBm���c��pso� !����s��e%�bS���
��JA��h� �����ﵰ���l }���D�Ģ����|zza)^���g�k�>�[z{fv��^���|إ�_����b��!�~Ɔ�zU�Uk�$R�^����L��֣�Y��;��N�\�p�o������R�l�S�
7|�^3�GܾY�s��������3P�.զ�7�]�SO��8DB��sG�A�>��j,/�,]��O��H�s���<���.4���&c�
���ż�!�'��̆y����7�%�	������ G�C�*[�IZ���z�#��ڡh�x=����=���'.!���.ύ�t�����ג�su3�e��̀�-�s9-TK)�6�$k�P3�۲F�� �����;D��F�B�wc�]�({�vz��� �K3�@�T��(��<�ۇH5�ORN�^5be�S����RpC�.l���P�8�²�)�kM�aS��Z��ԧ	��;�nF9�$�ϐP��e��hGZJ���藏:s���"�Ϩǔ�&2�Y����Sc~����'h��Wd{N��WnvB��V0qxNe�ŃQh�%�5��J[��N;K{��\Խ3
�I�����2aa� �����骓��sD�RIc6�>MK�sm5�isZܝ�H�G*!9�)(w�W���`vl������򏚡�*��o$���>D}�BC"1��a��if�2�#�9ܚ@OX)�ښOGĀX>��>ǘD���'b\�<�a#@���#�`�gv<�f]���pP4ܕK$���4��&ZQ(�w�B��0P�QC�J�(f\<kgj�����Q.0�LG�7�L�«��o��R�
(���HJ�����\3]�l���~���`��i���`��T%������"���=ΰ�����ե�����}�m:��8������G~ -�N��*� 1�cd[�/��A��
.,3���R	8����=/rW��a���@qc��	�Z0T[��w?�ʍ	�/+����oCO��Mh⏚E�!r
9d��R#��s ��rKk�hT�����O�t���y=F<��LOH$5+o�����3-��]�LE%?��7���k��E�]�rɃ��ժLj���X�hDP��U�z*臽> �λ4�lX���P�4��<��w�[�
���ɇ�@v[>���y�� �r:�
�j��hhk�2�՚ja|w?����9JUi$����S\�ͭ�h�}���@2���`���k+Δ��9E��pQ���#�t�ׅ�CJ�L++_@��R������B�n�j~h��N�yk,���<eԣ0�	���3�~�ڜΜk���iɘ8ȇ�:�Z�%Շ�9�r9(xO	�����'?�;|�\y�� �Ǣ�N��-��4�0F�����Ra)��Ʋ��<d��u��/��S�Wq�ڮ����>=<��C�kR	���X`����1��~�mk � ��M�ZT���F��}�8��ޤ�jb�x#�t2R��5
N����,��N��#U�&�W�������~@�V�Y�q�� }^_���gv3����:��Lt��c ���O*&�c��?떓	�v 9���vk{ؿF�]I����Jj�Y��0^��m⒡�覍\����E�p���k��8�hn�k$ig���ƓA�'��;��a��;oLZ�"�&��:,�W!N��B:�Y`�r�1%���g��-�N5�Kx�  �Lc��F.c����35l�����^��Ը�x�5%�yzĸ�o F��Fś��h�Pc��q�soA�?��<��J�|t#f�}i�����\sۆyE�>�W�ҧ\@�nI��յ�\�%1�N�����F-+?�B�������Q}�J��X9r�W���-ʇ�&������RݪwQŊmw��=p���G��=����n����)|gu ��_��M�wo��5�~��u���/(ڈ�qk���Чqi��1'�69��M�U���Ԍh�`��]��1	��TƧ4�OL�)��U�˥��X��Z2� a��eH��Q}X��-�VN��hǎ1h�$L�Lw�����l�=�8�ܒ��
;y
XXj��	�a�m=��#)��{�'g��#;��2&˨p1Ǹ*���6OO�P9~�\,fl�@�U!��!��8�a���q�}{|���O��F�rvd�"z��2����,��i�<�3�e�~7��~����zG�4Ǌ���iw���(mG�����T'5ˊ��q���4��q���{����|CR���G�	�+͓y�y/Q�8F��0&���a���Bf΂!�'L��g�
���>g�TK%�K�
�SꡅȐ�Շ�F>��.�6��R=��U�+_G�G��Q�BS	���jz��=�e�����q2��S4e�t��q��Z��8̓*������I=��ww
N��WK����F�A�G44+"3��/�E�iCQB�W����$��i�/��V��F�	UR��µ�$��-�ߜ����0��o;\� PV�f/�t7�8��+�)�`,Gn{�8�fgs|�`jbf/���:_d}X����*�z��k�9ih)��2d[�-H�c�d�R_C,	�Z���� H�������T�7r����Y�K��$��s�Vy�����	�ɭ?����_BcJ�Gi�Q8������y��̈��{]g��!�E�EU��ƛM�rS��2�|�T=s�����P�鲕Xz�8���=�e�%9�ĸ���f���ϸd�O�RN��t��Ԧ�|���W4{8<�о ��#drU��q���׀��+%(�aD�Ux�����L�OG|z/4ݕ��K�yǼ��K&(	4TY$1�"����S�SM~g��mWѡ=L�o0|?��E^�	��4��kn��<���p�&�P�c���`��<�BM��I���+}�=�_��:B��^�9�u�S3�&�e�h��e�͎��Q��D{�o�T"K3���i�a�[��s��G�-ZrG@���o�
:F�fs5�/D�"C|*���W�j"Gp���X�ECY��
��Y����L>
�B3g��������"RQ�@8|����k�q℃,���
��~.��n
Dcs"_o㾽d��]�:���V�8f��\,����B��zd^r��0wd�$�r�	f���� ��jҎ|�K�s3(P�
_v�L�-A�9�ZfSZ��5
Q���t���ZKdQ[_]�tu:7����<o�'�jB�[�@��<����-/�v:�,�K�l*й��f|�A�jΔ���De��9|vB}G����*��nU<�[W��k���t��6�o���n&z,��!3����bW�Z�2g��Q�,�<�5�N�2�����Nn$�(u(��.��D)���0_�2t�����/�d���Us�2o�PX���/�ޘ�8�~����9ܷ�A4�}jB���1L4���b�@����eu������5�9\U��N�䝺 &��ǗRnK��~�c��n��10���X\_�K�=�+tA�,�&��X�H�B�1��FȔ张�湰S�	ҙPP�$HQԐ8�'�X�����PX'9�f�!�n���7F���U�Qv5H �O����ݏ.(�Ȱ�4ݷ�^ͻҢ"����Jw�����"����ޕ+5M�&F��+z�x��Un��q��b��x�@i7rӀ���wM��/x�Kg�V��|�ߺi%s2�';��w��Ig�5�b��x���`�X;҅v���~6�]������䍆�z���ZxrΟ��Y	�J�C�|�/�E~t���Nr+ء�f�#���f��]��BHX��<H��0��?c ǡ�~[K�f�>�EzFSm��O�+��5�
�XxY�QwSy�ɭI�q�M�EtY��&���~�p���TX�0�������\�MaF��Ob�Bn���	c�����|�_@њ��de�����uM�i|�m3m�����L��J� D�+Ќ1��0; *��?��Oq�J�m�2�
Pb�'�A�e%W� Ir��i���֝l��QD"���l��� �)���a\F��q����8��1P�PMh�B��%�-~}�k<�,��$�����mJW�h